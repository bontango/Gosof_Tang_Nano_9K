--Copyright (C)2014-2025 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.11.01 (64-bit)
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9
--Device Version: C
--Created Time: Wed Apr  2 18:23:20 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_RAM16S is
    port (
        dout: out std_logic_vector(7 downto 0);
        wre: in std_logic;
        ad: in std_logic_vector(10 downto 0);
        di: in std_logic_vector(7 downto 0);
        clk: in std_logic
    );
end Gowin_RAM16S;

architecture Behavioral of Gowin_RAM16S is

    signal ad4_inv: std_logic;
    signal ad5_inv: std_logic;
    signal ad6_inv: std_logic;
    signal lut_f_0: std_logic;
    signal ad7_inv: std_logic;
    signal ad8_inv: std_logic;
    signal ad9_inv: std_logic;
    signal ad10_inv: std_logic;
    signal lut_f_1: std_logic;
    signal lut_f_2: std_logic;
    signal lut_f_3: std_logic;
    signal lut_f_4: std_logic;
    signal lut_f_5: std_logic;
    signal lut_f_6: std_logic;
    signal lut_f_7: std_logic;
    signal lut_f_8: std_logic;
    signal lut_f_9: std_logic;
    signal lut_f_10: std_logic;
    signal lut_f_11: std_logic;
    signal lut_f_12: std_logic;
    signal lut_f_13: std_logic;
    signal lut_f_14: std_logic;
    signal lut_f_15: std_logic;
    signal lut_f_16: std_logic;
    signal lut_f_17: std_logic;
    signal lut_f_18: std_logic;
    signal lut_f_19: std_logic;
    signal lut_f_20: std_logic;
    signal lut_f_21: std_logic;
    signal lut_f_22: std_logic;
    signal lut_f_23: std_logic;
    signal lut_f_24: std_logic;
    signal lut_f_25: std_logic;
    signal lut_f_26: std_logic;
    signal lut_f_27: std_logic;
    signal lut_f_28: std_logic;
    signal lut_f_29: std_logic;
    signal lut_f_30: std_logic;
    signal lut_f_31: std_logic;
    signal lut_f_32: std_logic;
    signal lut_f_33: std_logic;
    signal lut_f_34: std_logic;
    signal lut_f_35: std_logic;
    signal lut_f_36: std_logic;
    signal lut_f_37: std_logic;
    signal lut_f_38: std_logic;
    signal lut_f_39: std_logic;
    signal lut_f_40: std_logic;
    signal lut_f_41: std_logic;
    signal lut_f_42: std_logic;
    signal lut_f_43: std_logic;
    signal lut_f_44: std_logic;
    signal lut_f_45: std_logic;
    signal lut_f_46: std_logic;
    signal lut_f_47: std_logic;
    signal lut_f_48: std_logic;
    signal lut_f_49: std_logic;
    signal lut_f_50: std_logic;
    signal lut_f_51: std_logic;
    signal lut_f_52: std_logic;
    signal lut_f_53: std_logic;
    signal lut_f_54: std_logic;
    signal lut_f_55: std_logic;
    signal lut_f_56: std_logic;
    signal lut_f_57: std_logic;
    signal lut_f_58: std_logic;
    signal lut_f_59: std_logic;
    signal lut_f_60: std_logic;
    signal lut_f_61: std_logic;
    signal lut_f_62: std_logic;
    signal lut_f_63: std_logic;
    signal lut_f_64: std_logic;
    signal lut_f_65: std_logic;
    signal lut_f_66: std_logic;
    signal lut_f_67: std_logic;
    signal lut_f_68: std_logic;
    signal lut_f_69: std_logic;
    signal lut_f_70: std_logic;
    signal lut_f_71: std_logic;
    signal lut_f_72: std_logic;
    signal lut_f_73: std_logic;
    signal lut_f_74: std_logic;
    signal lut_f_75: std_logic;
    signal lut_f_76: std_logic;
    signal lut_f_77: std_logic;
    signal lut_f_78: std_logic;
    signal lut_f_79: std_logic;
    signal lut_f_80: std_logic;
    signal lut_f_81: std_logic;
    signal lut_f_82: std_logic;
    signal lut_f_83: std_logic;
    signal lut_f_84: std_logic;
    signal lut_f_85: std_logic;
    signal lut_f_86: std_logic;
    signal lut_f_87: std_logic;
    signal lut_f_88: std_logic;
    signal lut_f_89: std_logic;
    signal lut_f_90: std_logic;
    signal lut_f_91: std_logic;
    signal lut_f_92: std_logic;
    signal lut_f_93: std_logic;
    signal lut_f_94: std_logic;
    signal lut_f_95: std_logic;
    signal lut_f_96: std_logic;
    signal lut_f_97: std_logic;
    signal lut_f_98: std_logic;
    signal lut_f_99: std_logic;
    signal lut_f_100: std_logic;
    signal lut_f_101: std_logic;
    signal lut_f_102: std_logic;
    signal lut_f_103: std_logic;
    signal lut_f_104: std_logic;
    signal lut_f_105: std_logic;
    signal lut_f_106: std_logic;
    signal lut_f_107: std_logic;
    signal lut_f_108: std_logic;
    signal lut_f_109: std_logic;
    signal lut_f_110: std_logic;
    signal lut_f_111: std_logic;
    signal lut_f_112: std_logic;
    signal lut_f_113: std_logic;
    signal lut_f_114: std_logic;
    signal lut_f_115: std_logic;
    signal lut_f_116: std_logic;
    signal lut_f_117: std_logic;
    signal lut_f_118: std_logic;
    signal lut_f_119: std_logic;
    signal lut_f_120: std_logic;
    signal lut_f_121: std_logic;
    signal lut_f_122: std_logic;
    signal lut_f_123: std_logic;
    signal lut_f_124: std_logic;
    signal lut_f_125: std_logic;
    signal lut_f_126: std_logic;
    signal lut_f_127: std_logic;
    signal lut_f_128: std_logic;
    signal lut_f_129: std_logic;
    signal lut_f_130: std_logic;
    signal lut_f_131: std_logic;
    signal lut_f_132: std_logic;
    signal lut_f_133: std_logic;
    signal lut_f_134: std_logic;
    signal lut_f_135: std_logic;
    signal lut_f_136: std_logic;
    signal lut_f_137: std_logic;
    signal lut_f_138: std_logic;
    signal lut_f_139: std_logic;
    signal lut_f_140: std_logic;
    signal lut_f_141: std_logic;
    signal lut_f_142: std_logic;
    signal lut_f_143: std_logic;
    signal lut_f_144: std_logic;
    signal lut_f_145: std_logic;
    signal lut_f_146: std_logic;
    signal lut_f_147: std_logic;
    signal lut_f_148: std_logic;
    signal lut_f_149: std_logic;
    signal lut_f_150: std_logic;
    signal lut_f_151: std_logic;
    signal lut_f_152: std_logic;
    signal lut_f_153: std_logic;
    signal lut_f_154: std_logic;
    signal lut_f_155: std_logic;
    signal lut_f_156: std_logic;
    signal lut_f_157: std_logic;
    signal lut_f_158: std_logic;
    signal lut_f_159: std_logic;
    signal lut_f_160: std_logic;
    signal lut_f_161: std_logic;
    signal lut_f_162: std_logic;
    signal lut_f_163: std_logic;
    signal lut_f_164: std_logic;
    signal lut_f_165: std_logic;
    signal lut_f_166: std_logic;
    signal lut_f_167: std_logic;
    signal lut_f_168: std_logic;
    signal lut_f_169: std_logic;
    signal lut_f_170: std_logic;
    signal lut_f_171: std_logic;
    signal lut_f_172: std_logic;
    signal lut_f_173: std_logic;
    signal lut_f_174: std_logic;
    signal lut_f_175: std_logic;
    signal lut_f_176: std_logic;
    signal lut_f_177: std_logic;
    signal lut_f_178: std_logic;
    signal lut_f_179: std_logic;
    signal lut_f_180: std_logic;
    signal lut_f_181: std_logic;
    signal lut_f_182: std_logic;
    signal lut_f_183: std_logic;
    signal lut_f_184: std_logic;
    signal lut_f_185: std_logic;
    signal lut_f_186: std_logic;
    signal lut_f_187: std_logic;
    signal lut_f_188: std_logic;
    signal lut_f_189: std_logic;
    signal lut_f_190: std_logic;
    signal lut_f_191: std_logic;
    signal lut_f_192: std_logic;
    signal lut_f_193: std_logic;
    signal lut_f_194: std_logic;
    signal lut_f_195: std_logic;
    signal lut_f_196: std_logic;
    signal lut_f_197: std_logic;
    signal lut_f_198: std_logic;
    signal lut_f_199: std_logic;
    signal lut_f_200: std_logic;
    signal lut_f_201: std_logic;
    signal lut_f_202: std_logic;
    signal lut_f_203: std_logic;
    signal lut_f_204: std_logic;
    signal lut_f_205: std_logic;
    signal lut_f_206: std_logic;
    signal lut_f_207: std_logic;
    signal lut_f_208: std_logic;
    signal lut_f_209: std_logic;
    signal lut_f_210: std_logic;
    signal lut_f_211: std_logic;
    signal lut_f_212: std_logic;
    signal lut_f_213: std_logic;
    signal lut_f_214: std_logic;
    signal lut_f_215: std_logic;
    signal lut_f_216: std_logic;
    signal lut_f_217: std_logic;
    signal lut_f_218: std_logic;
    signal lut_f_219: std_logic;
    signal lut_f_220: std_logic;
    signal lut_f_221: std_logic;
    signal lut_f_222: std_logic;
    signal lut_f_223: std_logic;
    signal lut_f_224: std_logic;
    signal lut_f_225: std_logic;
    signal lut_f_226: std_logic;
    signal lut_f_227: std_logic;
    signal lut_f_228: std_logic;
    signal lut_f_229: std_logic;
    signal lut_f_230: std_logic;
    signal lut_f_231: std_logic;
    signal lut_f_232: std_logic;
    signal lut_f_233: std_logic;
    signal lut_f_234: std_logic;
    signal lut_f_235: std_logic;
    signal lut_f_236: std_logic;
    signal lut_f_237: std_logic;
    signal lut_f_238: std_logic;
    signal lut_f_239: std_logic;
    signal lut_f_240: std_logic;
    signal lut_f_241: std_logic;
    signal lut_f_242: std_logic;
    signal lut_f_243: std_logic;
    signal lut_f_244: std_logic;
    signal lut_f_245: std_logic;
    signal lut_f_246: std_logic;
    signal lut_f_247: std_logic;
    signal lut_f_248: std_logic;
    signal lut_f_249: std_logic;
    signal lut_f_250: std_logic;
    signal lut_f_251: std_logic;
    signal lut_f_252: std_logic;
    signal lut_f_253: std_logic;
    signal lut_f_254: std_logic;
    signal lut_f_255: std_logic;
    signal lut_f_256: std_logic;
    signal lut_f_257: std_logic;
    signal lut_f_258: std_logic;
    signal lut_f_259: std_logic;
    signal lut_f_260: std_logic;
    signal lut_f_261: std_logic;
    signal lut_f_262: std_logic;
    signal lut_f_263: std_logic;
    signal lut_f_264: std_logic;
    signal lut_f_265: std_logic;
    signal lut_f_266: std_logic;
    signal lut_f_267: std_logic;
    signal lut_f_268: std_logic;
    signal lut_f_269: std_logic;
    signal lut_f_270: std_logic;
    signal lut_f_271: std_logic;
    signal lut_f_272: std_logic;
    signal lut_f_273: std_logic;
    signal lut_f_274: std_logic;
    signal lut_f_275: std_logic;
    signal lut_f_276: std_logic;
    signal lut_f_277: std_logic;
    signal lut_f_278: std_logic;
    signal lut_f_279: std_logic;
    signal lut_f_280: std_logic;
    signal lut_f_281: std_logic;
    signal lut_f_282: std_logic;
    signal lut_f_283: std_logic;
    signal lut_f_284: std_logic;
    signal lut_f_285: std_logic;
    signal lut_f_286: std_logic;
    signal lut_f_287: std_logic;
    signal lut_f_288: std_logic;
    signal lut_f_289: std_logic;
    signal lut_f_290: std_logic;
    signal lut_f_291: std_logic;
    signal lut_f_292: std_logic;
    signal lut_f_293: std_logic;
    signal lut_f_294: std_logic;
    signal lut_f_295: std_logic;
    signal lut_f_296: std_logic;
    signal lut_f_297: std_logic;
    signal lut_f_298: std_logic;
    signal lut_f_299: std_logic;
    signal lut_f_300: std_logic;
    signal lut_f_301: std_logic;
    signal lut_f_302: std_logic;
    signal lut_f_303: std_logic;
    signal lut_f_304: std_logic;
    signal lut_f_305: std_logic;
    signal lut_f_306: std_logic;
    signal lut_f_307: std_logic;
    signal lut_f_308: std_logic;
    signal lut_f_309: std_logic;
    signal lut_f_310: std_logic;
    signal lut_f_311: std_logic;
    signal lut_f_312: std_logic;
    signal lut_f_313: std_logic;
    signal lut_f_314: std_logic;
    signal lut_f_315: std_logic;
    signal lut_f_316: std_logic;
    signal lut_f_317: std_logic;
    signal lut_f_318: std_logic;
    signal lut_f_319: std_logic;
    signal lut_f_320: std_logic;
    signal lut_f_321: std_logic;
    signal lut_f_322: std_logic;
    signal lut_f_323: std_logic;
    signal lut_f_324: std_logic;
    signal lut_f_325: std_logic;
    signal lut_f_326: std_logic;
    signal lut_f_327: std_logic;
    signal lut_f_328: std_logic;
    signal lut_f_329: std_logic;
    signal lut_f_330: std_logic;
    signal lut_f_331: std_logic;
    signal lut_f_332: std_logic;
    signal lut_f_333: std_logic;
    signal lut_f_334: std_logic;
    signal lut_f_335: std_logic;
    signal lut_f_336: std_logic;
    signal lut_f_337: std_logic;
    signal lut_f_338: std_logic;
    signal lut_f_339: std_logic;
    signal lut_f_340: std_logic;
    signal lut_f_341: std_logic;
    signal lut_f_342: std_logic;
    signal lut_f_343: std_logic;
    signal lut_f_344: std_logic;
    signal lut_f_345: std_logic;
    signal lut_f_346: std_logic;
    signal lut_f_347: std_logic;
    signal lut_f_348: std_logic;
    signal lut_f_349: std_logic;
    signal lut_f_350: std_logic;
    signal lut_f_351: std_logic;
    signal lut_f_352: std_logic;
    signal lut_f_353: std_logic;
    signal lut_f_354: std_logic;
    signal lut_f_355: std_logic;
    signal lut_f_356: std_logic;
    signal lut_f_357: std_logic;
    signal lut_f_358: std_logic;
    signal lut_f_359: std_logic;
    signal lut_f_360: std_logic;
    signal lut_f_361: std_logic;
    signal lut_f_362: std_logic;
    signal lut_f_363: std_logic;
    signal lut_f_364: std_logic;
    signal lut_f_365: std_logic;
    signal lut_f_366: std_logic;
    signal lut_f_367: std_logic;
    signal lut_f_368: std_logic;
    signal lut_f_369: std_logic;
    signal lut_f_370: std_logic;
    signal lut_f_371: std_logic;
    signal lut_f_372: std_logic;
    signal lut_f_373: std_logic;
    signal lut_f_374: std_logic;
    signal lut_f_375: std_logic;
    signal lut_f_376: std_logic;
    signal lut_f_377: std_logic;
    signal lut_f_378: std_logic;
    signal lut_f_379: std_logic;
    signal lut_f_380: std_logic;
    signal lut_f_381: std_logic;
    signal lut_f_382: std_logic;
    signal lut_f_383: std_logic;
    signal ram16s_inst_0_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_1_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_2_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_3_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_4_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_5_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_6_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_7_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_8_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_9_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_10_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_11_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_12_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_13_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_14_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_15_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_16_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_17_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_18_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_19_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_20_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_21_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_22_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_23_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_24_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_25_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_26_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_27_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_28_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_29_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_30_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_31_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_32_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_33_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_34_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_35_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_36_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_37_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_38_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_39_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_40_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_41_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_42_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_43_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_44_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_45_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_46_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_47_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_48_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_49_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_50_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_51_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_52_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_53_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_54_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_55_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_56_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_57_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_58_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_59_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_60_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_61_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_62_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_63_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_64_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_65_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_66_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_67_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_68_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_69_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_70_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_71_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_72_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_73_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_74_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_75_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_76_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_77_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_78_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_79_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_80_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_81_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_82_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_83_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_84_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_85_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_86_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_87_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_88_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_89_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_90_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_91_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_92_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_93_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_94_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_95_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_96_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_97_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_98_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_99_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_100_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_101_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_102_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_103_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_104_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_105_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_106_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_107_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_108_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_109_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_110_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_111_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_112_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_113_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_114_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_115_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_116_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_117_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_118_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_119_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_120_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_121_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_122_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_123_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_124_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_125_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_126_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_127_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_128_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_129_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_130_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_131_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_132_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_133_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_134_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_135_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_136_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_137_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_138_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_139_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_140_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_141_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_142_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_143_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_144_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_145_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_146_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_147_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_148_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_149_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_150_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_151_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_152_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_153_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_154_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_155_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_156_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_157_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_158_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_159_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_160_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_161_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_162_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_163_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_164_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_165_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_166_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_167_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_168_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_169_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_170_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_171_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_172_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_173_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_174_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_175_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_176_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_177_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_178_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_179_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_180_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_181_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_182_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_183_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_184_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_185_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_186_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_187_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_188_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_189_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_190_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_191_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_192_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_193_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_194_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_195_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_196_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_197_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_198_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_199_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_200_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_201_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_202_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_203_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_204_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_205_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_206_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_207_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_208_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_209_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_210_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_211_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_212_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_213_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_214_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_215_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_216_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_217_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_218_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_219_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_220_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_221_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_222_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_223_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_224_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_225_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_226_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_227_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_228_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_229_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_230_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_231_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_232_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_233_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_234_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_235_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_236_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_237_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_238_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_239_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_240_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_241_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_242_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_243_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_244_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_245_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_246_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_247_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_248_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_249_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_250_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_251_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_252_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_253_dout: std_logic_vector(7 downto 4);
    signal ram16s_inst_254_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_255_dout: std_logic_vector(7 downto 4);
    signal mux_o_0: std_logic;
    signal mux_o_1: std_logic;
    signal mux_o_2: std_logic;
    signal mux_o_3: std_logic;
    signal mux_o_4: std_logic;
    signal mux_o_5: std_logic;
    signal mux_o_6: std_logic;
    signal mux_o_7: std_logic;
    signal mux_o_8: std_logic;
    signal mux_o_9: std_logic;
    signal mux_o_10: std_logic;
    signal mux_o_11: std_logic;
    signal mux_o_12: std_logic;
    signal mux_o_13: std_logic;
    signal mux_o_14: std_logic;
    signal mux_o_15: std_logic;
    signal mux_o_16: std_logic;
    signal mux_o_17: std_logic;
    signal mux_o_18: std_logic;
    signal mux_o_19: std_logic;
    signal mux_o_20: std_logic;
    signal mux_o_21: std_logic;
    signal mux_o_22: std_logic;
    signal mux_o_23: std_logic;
    signal mux_o_24: std_logic;
    signal mux_o_25: std_logic;
    signal mux_o_26: std_logic;
    signal mux_o_27: std_logic;
    signal mux_o_28: std_logic;
    signal mux_o_29: std_logic;
    signal mux_o_30: std_logic;
    signal mux_o_31: std_logic;
    signal mux_o_32: std_logic;
    signal mux_o_33: std_logic;
    signal mux_o_34: std_logic;
    signal mux_o_35: std_logic;
    signal mux_o_36: std_logic;
    signal mux_o_37: std_logic;
    signal mux_o_38: std_logic;
    signal mux_o_39: std_logic;
    signal mux_o_40: std_logic;
    signal mux_o_41: std_logic;
    signal mux_o_42: std_logic;
    signal mux_o_43: std_logic;
    signal mux_o_44: std_logic;
    signal mux_o_45: std_logic;
    signal mux_o_46: std_logic;
    signal mux_o_47: std_logic;
    signal mux_o_48: std_logic;
    signal mux_o_49: std_logic;
    signal mux_o_50: std_logic;
    signal mux_o_51: std_logic;
    signal mux_o_52: std_logic;
    signal mux_o_53: std_logic;
    signal mux_o_54: std_logic;
    signal mux_o_55: std_logic;
    signal mux_o_56: std_logic;
    signal mux_o_57: std_logic;
    signal mux_o_58: std_logic;
    signal mux_o_59: std_logic;
    signal mux_o_60: std_logic;
    signal mux_o_61: std_logic;
    signal mux_o_62: std_logic;
    signal mux_o_63: std_logic;
    signal mux_o_64: std_logic;
    signal mux_o_65: std_logic;
    signal mux_o_66: std_logic;
    signal mux_o_67: std_logic;
    signal mux_o_68: std_logic;
    signal mux_o_69: std_logic;
    signal mux_o_70: std_logic;
    signal mux_o_71: std_logic;
    signal mux_o_72: std_logic;
    signal mux_o_73: std_logic;
    signal mux_o_74: std_logic;
    signal mux_o_75: std_logic;
    signal mux_o_76: std_logic;
    signal mux_o_77: std_logic;
    signal mux_o_78: std_logic;
    signal mux_o_79: std_logic;
    signal mux_o_80: std_logic;
    signal mux_o_81: std_logic;
    signal mux_o_82: std_logic;
    signal mux_o_83: std_logic;
    signal mux_o_84: std_logic;
    signal mux_o_85: std_logic;
    signal mux_o_86: std_logic;
    signal mux_o_87: std_logic;
    signal mux_o_88: std_logic;
    signal mux_o_89: std_logic;
    signal mux_o_90: std_logic;
    signal mux_o_91: std_logic;
    signal mux_o_92: std_logic;
    signal mux_o_93: std_logic;
    signal mux_o_94: std_logic;
    signal mux_o_95: std_logic;
    signal mux_o_96: std_logic;
    signal mux_o_97: std_logic;
    signal mux_o_98: std_logic;
    signal mux_o_99: std_logic;
    signal mux_o_100: std_logic;
    signal mux_o_101: std_logic;
    signal mux_o_102: std_logic;
    signal mux_o_103: std_logic;
    signal mux_o_104: std_logic;
    signal mux_o_105: std_logic;
    signal mux_o_106: std_logic;
    signal mux_o_107: std_logic;
    signal mux_o_108: std_logic;
    signal mux_o_109: std_logic;
    signal mux_o_110: std_logic;
    signal mux_o_111: std_logic;
    signal mux_o_112: std_logic;
    signal mux_o_113: std_logic;
    signal mux_o_114: std_logic;
    signal mux_o_115: std_logic;
    signal mux_o_116: std_logic;
    signal mux_o_117: std_logic;
    signal mux_o_118: std_logic;
    signal mux_o_119: std_logic;
    signal mux_o_120: std_logic;
    signal mux_o_121: std_logic;
    signal mux_o_122: std_logic;
    signal mux_o_123: std_logic;
    signal mux_o_124: std_logic;
    signal mux_o_125: std_logic;
    signal mux_o_127: std_logic;
    signal mux_o_128: std_logic;
    signal mux_o_129: std_logic;
    signal mux_o_130: std_logic;
    signal mux_o_131: std_logic;
    signal mux_o_132: std_logic;
    signal mux_o_133: std_logic;
    signal mux_o_134: std_logic;
    signal mux_o_135: std_logic;
    signal mux_o_136: std_logic;
    signal mux_o_137: std_logic;
    signal mux_o_138: std_logic;
    signal mux_o_139: std_logic;
    signal mux_o_140: std_logic;
    signal mux_o_141: std_logic;
    signal mux_o_142: std_logic;
    signal mux_o_143: std_logic;
    signal mux_o_144: std_logic;
    signal mux_o_145: std_logic;
    signal mux_o_146: std_logic;
    signal mux_o_147: std_logic;
    signal mux_o_148: std_logic;
    signal mux_o_149: std_logic;
    signal mux_o_150: std_logic;
    signal mux_o_151: std_logic;
    signal mux_o_152: std_logic;
    signal mux_o_153: std_logic;
    signal mux_o_154: std_logic;
    signal mux_o_155: std_logic;
    signal mux_o_156: std_logic;
    signal mux_o_157: std_logic;
    signal mux_o_158: std_logic;
    signal mux_o_159: std_logic;
    signal mux_o_160: std_logic;
    signal mux_o_161: std_logic;
    signal mux_o_162: std_logic;
    signal mux_o_163: std_logic;
    signal mux_o_164: std_logic;
    signal mux_o_165: std_logic;
    signal mux_o_166: std_logic;
    signal mux_o_167: std_logic;
    signal mux_o_168: std_logic;
    signal mux_o_169: std_logic;
    signal mux_o_170: std_logic;
    signal mux_o_171: std_logic;
    signal mux_o_172: std_logic;
    signal mux_o_173: std_logic;
    signal mux_o_174: std_logic;
    signal mux_o_175: std_logic;
    signal mux_o_176: std_logic;
    signal mux_o_177: std_logic;
    signal mux_o_178: std_logic;
    signal mux_o_179: std_logic;
    signal mux_o_180: std_logic;
    signal mux_o_181: std_logic;
    signal mux_o_182: std_logic;
    signal mux_o_183: std_logic;
    signal mux_o_184: std_logic;
    signal mux_o_185: std_logic;
    signal mux_o_186: std_logic;
    signal mux_o_187: std_logic;
    signal mux_o_188: std_logic;
    signal mux_o_189: std_logic;
    signal mux_o_190: std_logic;
    signal mux_o_191: std_logic;
    signal mux_o_192: std_logic;
    signal mux_o_193: std_logic;
    signal mux_o_194: std_logic;
    signal mux_o_195: std_logic;
    signal mux_o_196: std_logic;
    signal mux_o_197: std_logic;
    signal mux_o_198: std_logic;
    signal mux_o_199: std_logic;
    signal mux_o_200: std_logic;
    signal mux_o_201: std_logic;
    signal mux_o_202: std_logic;
    signal mux_o_203: std_logic;
    signal mux_o_204: std_logic;
    signal mux_o_205: std_logic;
    signal mux_o_206: std_logic;
    signal mux_o_207: std_logic;
    signal mux_o_208: std_logic;
    signal mux_o_209: std_logic;
    signal mux_o_210: std_logic;
    signal mux_o_211: std_logic;
    signal mux_o_212: std_logic;
    signal mux_o_213: std_logic;
    signal mux_o_214: std_logic;
    signal mux_o_215: std_logic;
    signal mux_o_216: std_logic;
    signal mux_o_217: std_logic;
    signal mux_o_218: std_logic;
    signal mux_o_219: std_logic;
    signal mux_o_220: std_logic;
    signal mux_o_221: std_logic;
    signal mux_o_222: std_logic;
    signal mux_o_223: std_logic;
    signal mux_o_224: std_logic;
    signal mux_o_225: std_logic;
    signal mux_o_226: std_logic;
    signal mux_o_227: std_logic;
    signal mux_o_228: std_logic;
    signal mux_o_229: std_logic;
    signal mux_o_230: std_logic;
    signal mux_o_231: std_logic;
    signal mux_o_232: std_logic;
    signal mux_o_233: std_logic;
    signal mux_o_234: std_logic;
    signal mux_o_235: std_logic;
    signal mux_o_236: std_logic;
    signal mux_o_237: std_logic;
    signal mux_o_238: std_logic;
    signal mux_o_239: std_logic;
    signal mux_o_240: std_logic;
    signal mux_o_241: std_logic;
    signal mux_o_242: std_logic;
    signal mux_o_243: std_logic;
    signal mux_o_244: std_logic;
    signal mux_o_245: std_logic;
    signal mux_o_246: std_logic;
    signal mux_o_247: std_logic;
    signal mux_o_248: std_logic;
    signal mux_o_249: std_logic;
    signal mux_o_250: std_logic;
    signal mux_o_251: std_logic;
    signal mux_o_252: std_logic;
    signal mux_o_254: std_logic;
    signal mux_o_255: std_logic;
    signal mux_o_256: std_logic;
    signal mux_o_257: std_logic;
    signal mux_o_258: std_logic;
    signal mux_o_259: std_logic;
    signal mux_o_260: std_logic;
    signal mux_o_261: std_logic;
    signal mux_o_262: std_logic;
    signal mux_o_263: std_logic;
    signal mux_o_264: std_logic;
    signal mux_o_265: std_logic;
    signal mux_o_266: std_logic;
    signal mux_o_267: std_logic;
    signal mux_o_268: std_logic;
    signal mux_o_269: std_logic;
    signal mux_o_270: std_logic;
    signal mux_o_271: std_logic;
    signal mux_o_272: std_logic;
    signal mux_o_273: std_logic;
    signal mux_o_274: std_logic;
    signal mux_o_275: std_logic;
    signal mux_o_276: std_logic;
    signal mux_o_277: std_logic;
    signal mux_o_278: std_logic;
    signal mux_o_279: std_logic;
    signal mux_o_280: std_logic;
    signal mux_o_281: std_logic;
    signal mux_o_282: std_logic;
    signal mux_o_283: std_logic;
    signal mux_o_284: std_logic;
    signal mux_o_285: std_logic;
    signal mux_o_286: std_logic;
    signal mux_o_287: std_logic;
    signal mux_o_288: std_logic;
    signal mux_o_289: std_logic;
    signal mux_o_290: std_logic;
    signal mux_o_291: std_logic;
    signal mux_o_292: std_logic;
    signal mux_o_293: std_logic;
    signal mux_o_294: std_logic;
    signal mux_o_295: std_logic;
    signal mux_o_296: std_logic;
    signal mux_o_297: std_logic;
    signal mux_o_298: std_logic;
    signal mux_o_299: std_logic;
    signal mux_o_300: std_logic;
    signal mux_o_301: std_logic;
    signal mux_o_302: std_logic;
    signal mux_o_303: std_logic;
    signal mux_o_304: std_logic;
    signal mux_o_305: std_logic;
    signal mux_o_306: std_logic;
    signal mux_o_307: std_logic;
    signal mux_o_308: std_logic;
    signal mux_o_309: std_logic;
    signal mux_o_310: std_logic;
    signal mux_o_311: std_logic;
    signal mux_o_312: std_logic;
    signal mux_o_313: std_logic;
    signal mux_o_314: std_logic;
    signal mux_o_315: std_logic;
    signal mux_o_316: std_logic;
    signal mux_o_317: std_logic;
    signal mux_o_318: std_logic;
    signal mux_o_319: std_logic;
    signal mux_o_320: std_logic;
    signal mux_o_321: std_logic;
    signal mux_o_322: std_logic;
    signal mux_o_323: std_logic;
    signal mux_o_324: std_logic;
    signal mux_o_325: std_logic;
    signal mux_o_326: std_logic;
    signal mux_o_327: std_logic;
    signal mux_o_328: std_logic;
    signal mux_o_329: std_logic;
    signal mux_o_330: std_logic;
    signal mux_o_331: std_logic;
    signal mux_o_332: std_logic;
    signal mux_o_333: std_logic;
    signal mux_o_334: std_logic;
    signal mux_o_335: std_logic;
    signal mux_o_336: std_logic;
    signal mux_o_337: std_logic;
    signal mux_o_338: std_logic;
    signal mux_o_339: std_logic;
    signal mux_o_340: std_logic;
    signal mux_o_341: std_logic;
    signal mux_o_342: std_logic;
    signal mux_o_343: std_logic;
    signal mux_o_344: std_logic;
    signal mux_o_345: std_logic;
    signal mux_o_346: std_logic;
    signal mux_o_347: std_logic;
    signal mux_o_348: std_logic;
    signal mux_o_349: std_logic;
    signal mux_o_350: std_logic;
    signal mux_o_351: std_logic;
    signal mux_o_352: std_logic;
    signal mux_o_353: std_logic;
    signal mux_o_354: std_logic;
    signal mux_o_355: std_logic;
    signal mux_o_356: std_logic;
    signal mux_o_357: std_logic;
    signal mux_o_358: std_logic;
    signal mux_o_359: std_logic;
    signal mux_o_360: std_logic;
    signal mux_o_361: std_logic;
    signal mux_o_362: std_logic;
    signal mux_o_363: std_logic;
    signal mux_o_364: std_logic;
    signal mux_o_365: std_logic;
    signal mux_o_366: std_logic;
    signal mux_o_367: std_logic;
    signal mux_o_368: std_logic;
    signal mux_o_369: std_logic;
    signal mux_o_370: std_logic;
    signal mux_o_371: std_logic;
    signal mux_o_372: std_logic;
    signal mux_o_373: std_logic;
    signal mux_o_374: std_logic;
    signal mux_o_375: std_logic;
    signal mux_o_376: std_logic;
    signal mux_o_377: std_logic;
    signal mux_o_378: std_logic;
    signal mux_o_379: std_logic;
    signal mux_o_381: std_logic;
    signal mux_o_382: std_logic;
    signal mux_o_383: std_logic;
    signal mux_o_384: std_logic;
    signal mux_o_385: std_logic;
    signal mux_o_386: std_logic;
    signal mux_o_387: std_logic;
    signal mux_o_388: std_logic;
    signal mux_o_389: std_logic;
    signal mux_o_390: std_logic;
    signal mux_o_391: std_logic;
    signal mux_o_392: std_logic;
    signal mux_o_393: std_logic;
    signal mux_o_394: std_logic;
    signal mux_o_395: std_logic;
    signal mux_o_396: std_logic;
    signal mux_o_397: std_logic;
    signal mux_o_398: std_logic;
    signal mux_o_399: std_logic;
    signal mux_o_400: std_logic;
    signal mux_o_401: std_logic;
    signal mux_o_402: std_logic;
    signal mux_o_403: std_logic;
    signal mux_o_404: std_logic;
    signal mux_o_405: std_logic;
    signal mux_o_406: std_logic;
    signal mux_o_407: std_logic;
    signal mux_o_408: std_logic;
    signal mux_o_409: std_logic;
    signal mux_o_410: std_logic;
    signal mux_o_411: std_logic;
    signal mux_o_412: std_logic;
    signal mux_o_413: std_logic;
    signal mux_o_414: std_logic;
    signal mux_o_415: std_logic;
    signal mux_o_416: std_logic;
    signal mux_o_417: std_logic;
    signal mux_o_418: std_logic;
    signal mux_o_419: std_logic;
    signal mux_o_420: std_logic;
    signal mux_o_421: std_logic;
    signal mux_o_422: std_logic;
    signal mux_o_423: std_logic;
    signal mux_o_424: std_logic;
    signal mux_o_425: std_logic;
    signal mux_o_426: std_logic;
    signal mux_o_427: std_logic;
    signal mux_o_428: std_logic;
    signal mux_o_429: std_logic;
    signal mux_o_430: std_logic;
    signal mux_o_431: std_logic;
    signal mux_o_432: std_logic;
    signal mux_o_433: std_logic;
    signal mux_o_434: std_logic;
    signal mux_o_435: std_logic;
    signal mux_o_436: std_logic;
    signal mux_o_437: std_logic;
    signal mux_o_438: std_logic;
    signal mux_o_439: std_logic;
    signal mux_o_440: std_logic;
    signal mux_o_441: std_logic;
    signal mux_o_442: std_logic;
    signal mux_o_443: std_logic;
    signal mux_o_444: std_logic;
    signal mux_o_445: std_logic;
    signal mux_o_446: std_logic;
    signal mux_o_447: std_logic;
    signal mux_o_448: std_logic;
    signal mux_o_449: std_logic;
    signal mux_o_450: std_logic;
    signal mux_o_451: std_logic;
    signal mux_o_452: std_logic;
    signal mux_o_453: std_logic;
    signal mux_o_454: std_logic;
    signal mux_o_455: std_logic;
    signal mux_o_456: std_logic;
    signal mux_o_457: std_logic;
    signal mux_o_458: std_logic;
    signal mux_o_459: std_logic;
    signal mux_o_460: std_logic;
    signal mux_o_461: std_logic;
    signal mux_o_462: std_logic;
    signal mux_o_463: std_logic;
    signal mux_o_464: std_logic;
    signal mux_o_465: std_logic;
    signal mux_o_466: std_logic;
    signal mux_o_467: std_logic;
    signal mux_o_468: std_logic;
    signal mux_o_469: std_logic;
    signal mux_o_470: std_logic;
    signal mux_o_471: std_logic;
    signal mux_o_472: std_logic;
    signal mux_o_473: std_logic;
    signal mux_o_474: std_logic;
    signal mux_o_475: std_logic;
    signal mux_o_476: std_logic;
    signal mux_o_477: std_logic;
    signal mux_o_478: std_logic;
    signal mux_o_479: std_logic;
    signal mux_o_480: std_logic;
    signal mux_o_481: std_logic;
    signal mux_o_482: std_logic;
    signal mux_o_483: std_logic;
    signal mux_o_484: std_logic;
    signal mux_o_485: std_logic;
    signal mux_o_486: std_logic;
    signal mux_o_487: std_logic;
    signal mux_o_488: std_logic;
    signal mux_o_489: std_logic;
    signal mux_o_490: std_logic;
    signal mux_o_491: std_logic;
    signal mux_o_492: std_logic;
    signal mux_o_493: std_logic;
    signal mux_o_494: std_logic;
    signal mux_o_495: std_logic;
    signal mux_o_496: std_logic;
    signal mux_o_497: std_logic;
    signal mux_o_498: std_logic;
    signal mux_o_499: std_logic;
    signal mux_o_500: std_logic;
    signal mux_o_501: std_logic;
    signal mux_o_502: std_logic;
    signal mux_o_503: std_logic;
    signal mux_o_504: std_logic;
    signal mux_o_505: std_logic;
    signal mux_o_506: std_logic;
    signal mux_o_508: std_logic;
    signal mux_o_509: std_logic;
    signal mux_o_510: std_logic;
    signal mux_o_511: std_logic;
    signal mux_o_512: std_logic;
    signal mux_o_513: std_logic;
    signal mux_o_514: std_logic;
    signal mux_o_515: std_logic;
    signal mux_o_516: std_logic;
    signal mux_o_517: std_logic;
    signal mux_o_518: std_logic;
    signal mux_o_519: std_logic;
    signal mux_o_520: std_logic;
    signal mux_o_521: std_logic;
    signal mux_o_522: std_logic;
    signal mux_o_523: std_logic;
    signal mux_o_524: std_logic;
    signal mux_o_525: std_logic;
    signal mux_o_526: std_logic;
    signal mux_o_527: std_logic;
    signal mux_o_528: std_logic;
    signal mux_o_529: std_logic;
    signal mux_o_530: std_logic;
    signal mux_o_531: std_logic;
    signal mux_o_532: std_logic;
    signal mux_o_533: std_logic;
    signal mux_o_534: std_logic;
    signal mux_o_535: std_logic;
    signal mux_o_536: std_logic;
    signal mux_o_537: std_logic;
    signal mux_o_538: std_logic;
    signal mux_o_539: std_logic;
    signal mux_o_540: std_logic;
    signal mux_o_541: std_logic;
    signal mux_o_542: std_logic;
    signal mux_o_543: std_logic;
    signal mux_o_544: std_logic;
    signal mux_o_545: std_logic;
    signal mux_o_546: std_logic;
    signal mux_o_547: std_logic;
    signal mux_o_548: std_logic;
    signal mux_o_549: std_logic;
    signal mux_o_550: std_logic;
    signal mux_o_551: std_logic;
    signal mux_o_552: std_logic;
    signal mux_o_553: std_logic;
    signal mux_o_554: std_logic;
    signal mux_o_555: std_logic;
    signal mux_o_556: std_logic;
    signal mux_o_557: std_logic;
    signal mux_o_558: std_logic;
    signal mux_o_559: std_logic;
    signal mux_o_560: std_logic;
    signal mux_o_561: std_logic;
    signal mux_o_562: std_logic;
    signal mux_o_563: std_logic;
    signal mux_o_564: std_logic;
    signal mux_o_565: std_logic;
    signal mux_o_566: std_logic;
    signal mux_o_567: std_logic;
    signal mux_o_568: std_logic;
    signal mux_o_569: std_logic;
    signal mux_o_570: std_logic;
    signal mux_o_571: std_logic;
    signal mux_o_572: std_logic;
    signal mux_o_573: std_logic;
    signal mux_o_574: std_logic;
    signal mux_o_575: std_logic;
    signal mux_o_576: std_logic;
    signal mux_o_577: std_logic;
    signal mux_o_578: std_logic;
    signal mux_o_579: std_logic;
    signal mux_o_580: std_logic;
    signal mux_o_581: std_logic;
    signal mux_o_582: std_logic;
    signal mux_o_583: std_logic;
    signal mux_o_584: std_logic;
    signal mux_o_585: std_logic;
    signal mux_o_586: std_logic;
    signal mux_o_587: std_logic;
    signal mux_o_588: std_logic;
    signal mux_o_589: std_logic;
    signal mux_o_590: std_logic;
    signal mux_o_591: std_logic;
    signal mux_o_592: std_logic;
    signal mux_o_593: std_logic;
    signal mux_o_594: std_logic;
    signal mux_o_595: std_logic;
    signal mux_o_596: std_logic;
    signal mux_o_597: std_logic;
    signal mux_o_598: std_logic;
    signal mux_o_599: std_logic;
    signal mux_o_600: std_logic;
    signal mux_o_601: std_logic;
    signal mux_o_602: std_logic;
    signal mux_o_603: std_logic;
    signal mux_o_604: std_logic;
    signal mux_o_605: std_logic;
    signal mux_o_606: std_logic;
    signal mux_o_607: std_logic;
    signal mux_o_608: std_logic;
    signal mux_o_609: std_logic;
    signal mux_o_610: std_logic;
    signal mux_o_611: std_logic;
    signal mux_o_612: std_logic;
    signal mux_o_613: std_logic;
    signal mux_o_614: std_logic;
    signal mux_o_615: std_logic;
    signal mux_o_616: std_logic;
    signal mux_o_617: std_logic;
    signal mux_o_618: std_logic;
    signal mux_o_619: std_logic;
    signal mux_o_620: std_logic;
    signal mux_o_621: std_logic;
    signal mux_o_622: std_logic;
    signal mux_o_623: std_logic;
    signal mux_o_624: std_logic;
    signal mux_o_625: std_logic;
    signal mux_o_626: std_logic;
    signal mux_o_627: std_logic;
    signal mux_o_628: std_logic;
    signal mux_o_629: std_logic;
    signal mux_o_630: std_logic;
    signal mux_o_631: std_logic;
    signal mux_o_632: std_logic;
    signal mux_o_633: std_logic;
    signal mux_o_635: std_logic;
    signal mux_o_636: std_logic;
    signal mux_o_637: std_logic;
    signal mux_o_638: std_logic;
    signal mux_o_639: std_logic;
    signal mux_o_640: std_logic;
    signal mux_o_641: std_logic;
    signal mux_o_642: std_logic;
    signal mux_o_643: std_logic;
    signal mux_o_644: std_logic;
    signal mux_o_645: std_logic;
    signal mux_o_646: std_logic;
    signal mux_o_647: std_logic;
    signal mux_o_648: std_logic;
    signal mux_o_649: std_logic;
    signal mux_o_650: std_logic;
    signal mux_o_651: std_logic;
    signal mux_o_652: std_logic;
    signal mux_o_653: std_logic;
    signal mux_o_654: std_logic;
    signal mux_o_655: std_logic;
    signal mux_o_656: std_logic;
    signal mux_o_657: std_logic;
    signal mux_o_658: std_logic;
    signal mux_o_659: std_logic;
    signal mux_o_660: std_logic;
    signal mux_o_661: std_logic;
    signal mux_o_662: std_logic;
    signal mux_o_663: std_logic;
    signal mux_o_664: std_logic;
    signal mux_o_665: std_logic;
    signal mux_o_666: std_logic;
    signal mux_o_667: std_logic;
    signal mux_o_668: std_logic;
    signal mux_o_669: std_logic;
    signal mux_o_670: std_logic;
    signal mux_o_671: std_logic;
    signal mux_o_672: std_logic;
    signal mux_o_673: std_logic;
    signal mux_o_674: std_logic;
    signal mux_o_675: std_logic;
    signal mux_o_676: std_logic;
    signal mux_o_677: std_logic;
    signal mux_o_678: std_logic;
    signal mux_o_679: std_logic;
    signal mux_o_680: std_logic;
    signal mux_o_681: std_logic;
    signal mux_o_682: std_logic;
    signal mux_o_683: std_logic;
    signal mux_o_684: std_logic;
    signal mux_o_685: std_logic;
    signal mux_o_686: std_logic;
    signal mux_o_687: std_logic;
    signal mux_o_688: std_logic;
    signal mux_o_689: std_logic;
    signal mux_o_690: std_logic;
    signal mux_o_691: std_logic;
    signal mux_o_692: std_logic;
    signal mux_o_693: std_logic;
    signal mux_o_694: std_logic;
    signal mux_o_695: std_logic;
    signal mux_o_696: std_logic;
    signal mux_o_697: std_logic;
    signal mux_o_698: std_logic;
    signal mux_o_699: std_logic;
    signal mux_o_700: std_logic;
    signal mux_o_701: std_logic;
    signal mux_o_702: std_logic;
    signal mux_o_703: std_logic;
    signal mux_o_704: std_logic;
    signal mux_o_705: std_logic;
    signal mux_o_706: std_logic;
    signal mux_o_707: std_logic;
    signal mux_o_708: std_logic;
    signal mux_o_709: std_logic;
    signal mux_o_710: std_logic;
    signal mux_o_711: std_logic;
    signal mux_o_712: std_logic;
    signal mux_o_713: std_logic;
    signal mux_o_714: std_logic;
    signal mux_o_715: std_logic;
    signal mux_o_716: std_logic;
    signal mux_o_717: std_logic;
    signal mux_o_718: std_logic;
    signal mux_o_719: std_logic;
    signal mux_o_720: std_logic;
    signal mux_o_721: std_logic;
    signal mux_o_722: std_logic;
    signal mux_o_723: std_logic;
    signal mux_o_724: std_logic;
    signal mux_o_725: std_logic;
    signal mux_o_726: std_logic;
    signal mux_o_727: std_logic;
    signal mux_o_728: std_logic;
    signal mux_o_729: std_logic;
    signal mux_o_730: std_logic;
    signal mux_o_731: std_logic;
    signal mux_o_732: std_logic;
    signal mux_o_733: std_logic;
    signal mux_o_734: std_logic;
    signal mux_o_735: std_logic;
    signal mux_o_736: std_logic;
    signal mux_o_737: std_logic;
    signal mux_o_738: std_logic;
    signal mux_o_739: std_logic;
    signal mux_o_740: std_logic;
    signal mux_o_741: std_logic;
    signal mux_o_742: std_logic;
    signal mux_o_743: std_logic;
    signal mux_o_744: std_logic;
    signal mux_o_745: std_logic;
    signal mux_o_746: std_logic;
    signal mux_o_747: std_logic;
    signal mux_o_748: std_logic;
    signal mux_o_749: std_logic;
    signal mux_o_750: std_logic;
    signal mux_o_751: std_logic;
    signal mux_o_752: std_logic;
    signal mux_o_753: std_logic;
    signal mux_o_754: std_logic;
    signal mux_o_755: std_logic;
    signal mux_o_756: std_logic;
    signal mux_o_757: std_logic;
    signal mux_o_758: std_logic;
    signal mux_o_759: std_logic;
    signal mux_o_760: std_logic;
    signal mux_o_762: std_logic;
    signal mux_o_763: std_logic;
    signal mux_o_764: std_logic;
    signal mux_o_765: std_logic;
    signal mux_o_766: std_logic;
    signal mux_o_767: std_logic;
    signal mux_o_768: std_logic;
    signal mux_o_769: std_logic;
    signal mux_o_770: std_logic;
    signal mux_o_771: std_logic;
    signal mux_o_772: std_logic;
    signal mux_o_773: std_logic;
    signal mux_o_774: std_logic;
    signal mux_o_775: std_logic;
    signal mux_o_776: std_logic;
    signal mux_o_777: std_logic;
    signal mux_o_778: std_logic;
    signal mux_o_779: std_logic;
    signal mux_o_780: std_logic;
    signal mux_o_781: std_logic;
    signal mux_o_782: std_logic;
    signal mux_o_783: std_logic;
    signal mux_o_784: std_logic;
    signal mux_o_785: std_logic;
    signal mux_o_786: std_logic;
    signal mux_o_787: std_logic;
    signal mux_o_788: std_logic;
    signal mux_o_789: std_logic;
    signal mux_o_790: std_logic;
    signal mux_o_791: std_logic;
    signal mux_o_792: std_logic;
    signal mux_o_793: std_logic;
    signal mux_o_794: std_logic;
    signal mux_o_795: std_logic;
    signal mux_o_796: std_logic;
    signal mux_o_797: std_logic;
    signal mux_o_798: std_logic;
    signal mux_o_799: std_logic;
    signal mux_o_800: std_logic;
    signal mux_o_801: std_logic;
    signal mux_o_802: std_logic;
    signal mux_o_803: std_logic;
    signal mux_o_804: std_logic;
    signal mux_o_805: std_logic;
    signal mux_o_806: std_logic;
    signal mux_o_807: std_logic;
    signal mux_o_808: std_logic;
    signal mux_o_809: std_logic;
    signal mux_o_810: std_logic;
    signal mux_o_811: std_logic;
    signal mux_o_812: std_logic;
    signal mux_o_813: std_logic;
    signal mux_o_814: std_logic;
    signal mux_o_815: std_logic;
    signal mux_o_816: std_logic;
    signal mux_o_817: std_logic;
    signal mux_o_818: std_logic;
    signal mux_o_819: std_logic;
    signal mux_o_820: std_logic;
    signal mux_o_821: std_logic;
    signal mux_o_822: std_logic;
    signal mux_o_823: std_logic;
    signal mux_o_824: std_logic;
    signal mux_o_825: std_logic;
    signal mux_o_826: std_logic;
    signal mux_o_827: std_logic;
    signal mux_o_828: std_logic;
    signal mux_o_829: std_logic;
    signal mux_o_830: std_logic;
    signal mux_o_831: std_logic;
    signal mux_o_832: std_logic;
    signal mux_o_833: std_logic;
    signal mux_o_834: std_logic;
    signal mux_o_835: std_logic;
    signal mux_o_836: std_logic;
    signal mux_o_837: std_logic;
    signal mux_o_838: std_logic;
    signal mux_o_839: std_logic;
    signal mux_o_840: std_logic;
    signal mux_o_841: std_logic;
    signal mux_o_842: std_logic;
    signal mux_o_843: std_logic;
    signal mux_o_844: std_logic;
    signal mux_o_845: std_logic;
    signal mux_o_846: std_logic;
    signal mux_o_847: std_logic;
    signal mux_o_848: std_logic;
    signal mux_o_849: std_logic;
    signal mux_o_850: std_logic;
    signal mux_o_851: std_logic;
    signal mux_o_852: std_logic;
    signal mux_o_853: std_logic;
    signal mux_o_854: std_logic;
    signal mux_o_855: std_logic;
    signal mux_o_856: std_logic;
    signal mux_o_857: std_logic;
    signal mux_o_858: std_logic;
    signal mux_o_859: std_logic;
    signal mux_o_860: std_logic;
    signal mux_o_861: std_logic;
    signal mux_o_862: std_logic;
    signal mux_o_863: std_logic;
    signal mux_o_864: std_logic;
    signal mux_o_865: std_logic;
    signal mux_o_866: std_logic;
    signal mux_o_867: std_logic;
    signal mux_o_868: std_logic;
    signal mux_o_869: std_logic;
    signal mux_o_870: std_logic;
    signal mux_o_871: std_logic;
    signal mux_o_872: std_logic;
    signal mux_o_873: std_logic;
    signal mux_o_874: std_logic;
    signal mux_o_875: std_logic;
    signal mux_o_876: std_logic;
    signal mux_o_877: std_logic;
    signal mux_o_878: std_logic;
    signal mux_o_879: std_logic;
    signal mux_o_880: std_logic;
    signal mux_o_881: std_logic;
    signal mux_o_882: std_logic;
    signal mux_o_883: std_logic;
    signal mux_o_884: std_logic;
    signal mux_o_885: std_logic;
    signal mux_o_886: std_logic;
    signal mux_o_887: std_logic;
    signal mux_o_889: std_logic;
    signal mux_o_890: std_logic;
    signal mux_o_891: std_logic;
    signal mux_o_892: std_logic;
    signal mux_o_893: std_logic;
    signal mux_o_894: std_logic;
    signal mux_o_895: std_logic;
    signal mux_o_896: std_logic;
    signal mux_o_897: std_logic;
    signal mux_o_898: std_logic;
    signal mux_o_899: std_logic;
    signal mux_o_900: std_logic;
    signal mux_o_901: std_logic;
    signal mux_o_902: std_logic;
    signal mux_o_903: std_logic;
    signal mux_o_904: std_logic;
    signal mux_o_905: std_logic;
    signal mux_o_906: std_logic;
    signal mux_o_907: std_logic;
    signal mux_o_908: std_logic;
    signal mux_o_909: std_logic;
    signal mux_o_910: std_logic;
    signal mux_o_911: std_logic;
    signal mux_o_912: std_logic;
    signal mux_o_913: std_logic;
    signal mux_o_914: std_logic;
    signal mux_o_915: std_logic;
    signal mux_o_916: std_logic;
    signal mux_o_917: std_logic;
    signal mux_o_918: std_logic;
    signal mux_o_919: std_logic;
    signal mux_o_920: std_logic;
    signal mux_o_921: std_logic;
    signal mux_o_922: std_logic;
    signal mux_o_923: std_logic;
    signal mux_o_924: std_logic;
    signal mux_o_925: std_logic;
    signal mux_o_926: std_logic;
    signal mux_o_927: std_logic;
    signal mux_o_928: std_logic;
    signal mux_o_929: std_logic;
    signal mux_o_930: std_logic;
    signal mux_o_931: std_logic;
    signal mux_o_932: std_logic;
    signal mux_o_933: std_logic;
    signal mux_o_934: std_logic;
    signal mux_o_935: std_logic;
    signal mux_o_936: std_logic;
    signal mux_o_937: std_logic;
    signal mux_o_938: std_logic;
    signal mux_o_939: std_logic;
    signal mux_o_940: std_logic;
    signal mux_o_941: std_logic;
    signal mux_o_942: std_logic;
    signal mux_o_943: std_logic;
    signal mux_o_944: std_logic;
    signal mux_o_945: std_logic;
    signal mux_o_946: std_logic;
    signal mux_o_947: std_logic;
    signal mux_o_948: std_logic;
    signal mux_o_949: std_logic;
    signal mux_o_950: std_logic;
    signal mux_o_951: std_logic;
    signal mux_o_952: std_logic;
    signal mux_o_953: std_logic;
    signal mux_o_954: std_logic;
    signal mux_o_955: std_logic;
    signal mux_o_956: std_logic;
    signal mux_o_957: std_logic;
    signal mux_o_958: std_logic;
    signal mux_o_959: std_logic;
    signal mux_o_960: std_logic;
    signal mux_o_961: std_logic;
    signal mux_o_962: std_logic;
    signal mux_o_963: std_logic;
    signal mux_o_964: std_logic;
    signal mux_o_965: std_logic;
    signal mux_o_966: std_logic;
    signal mux_o_967: std_logic;
    signal mux_o_968: std_logic;
    signal mux_o_969: std_logic;
    signal mux_o_970: std_logic;
    signal mux_o_971: std_logic;
    signal mux_o_972: std_logic;
    signal mux_o_973: std_logic;
    signal mux_o_974: std_logic;
    signal mux_o_975: std_logic;
    signal mux_o_976: std_logic;
    signal mux_o_977: std_logic;
    signal mux_o_978: std_logic;
    signal mux_o_979: std_logic;
    signal mux_o_980: std_logic;
    signal mux_o_981: std_logic;
    signal mux_o_982: std_logic;
    signal mux_o_983: std_logic;
    signal mux_o_984: std_logic;
    signal mux_o_985: std_logic;
    signal mux_o_986: std_logic;
    signal mux_o_987: std_logic;
    signal mux_o_988: std_logic;
    signal mux_o_989: std_logic;
    signal mux_o_990: std_logic;
    signal mux_o_991: std_logic;
    signal mux_o_992: std_logic;
    signal mux_o_993: std_logic;
    signal mux_o_994: std_logic;
    signal mux_o_995: std_logic;
    signal mux_o_996: std_logic;
    signal mux_o_997: std_logic;
    signal mux_o_998: std_logic;
    signal mux_o_999: std_logic;
    signal mux_o_1000: std_logic;
    signal mux_o_1001: std_logic;
    signal mux_o_1002: std_logic;
    signal mux_o_1003: std_logic;
    signal mux_o_1004: std_logic;
    signal mux_o_1005: std_logic;
    signal mux_o_1006: std_logic;
    signal mux_o_1007: std_logic;
    signal mux_o_1008: std_logic;
    signal mux_o_1009: std_logic;
    signal mux_o_1010: std_logic;
    signal mux_o_1011: std_logic;
    signal mux_o_1012: std_logic;
    signal mux_o_1013: std_logic;
    signal mux_o_1014: std_logic;
    signal gw_vcc: std_logic;

    -- component declaration
    component INV
        port (I: in std_logic; O: out std_logic);
    end component;

    -- component declaration
    component LUT4
        generic (
            INIT: in bit_vector := X"0000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic
        );
    end component;

    --component declaration
    component RAM16S4
        GENERIC ( INIT_0 : bit_vector(15 downto 0) := X"0000";
                  INIT_1 : bit_vector(15 downto 0) := X"0000";
                  INIT_2 : bit_vector(15 downto 0) := X"0000";
                  INIT_3 : bit_vector(15 downto 0) := X"0000"
        );
        port (
            DO: out std_logic_vector(3 downto 0);
            DI: in std_logic_vector(3 downto 0);
            AD: in std_logic_vector(3 downto 0);
            WRE: in std_logic;
            CLK: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    gw_vcc <= '1';

    inv_inst_0 : INV
        port map (I => ad(4), O => ad4_inv);

    inv_inst_1 : INV
        port map (I => ad(5), O => ad5_inv);

    inv_inst_2 : INV
        port map (I => ad(6), O => ad6_inv);

    inv_inst_3 : INV
        port map (I => ad(7), O => ad7_inv);

    inv_inst_4 : INV
        port map (I => ad(8), O => ad8_inv);

    inv_inst_5 : INV
        port map (I => ad(9), O => ad9_inv);

    inv_inst_6 : INV
        port map (I => ad(10), O => ad10_inv);

    lut_inst_0 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_0,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_1 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_1,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_2 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_2,
            I0 => lut_f_0,
            I1 => lut_f_1,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_3 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_3,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_4 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_4,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_5 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_5,
            I0 => lut_f_3,
            I1 => lut_f_4,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_6 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_6,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_7 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_7,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_8 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_8,
            I0 => lut_f_6,
            I1 => lut_f_7,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_9 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_9,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_10 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_10,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_11 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_11,
            I0 => lut_f_9,
            I1 => lut_f_10,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_12 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_12,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_13 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_13,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_14 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_14,
            I0 => lut_f_12,
            I1 => lut_f_13,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_15 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_15,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_16 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_16,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_17 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_17,
            I0 => lut_f_15,
            I1 => lut_f_16,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_18 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_18,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_19 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_19,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_20 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_20,
            I0 => lut_f_18,
            I1 => lut_f_19,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_21 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_21,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_22 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_22,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_23 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_23,
            I0 => lut_f_21,
            I1 => lut_f_22,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_24 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_24,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_25 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_25,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_26 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_26,
            I0 => lut_f_24,
            I1 => lut_f_25,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_27 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_27,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_28 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_28,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_29 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_29,
            I0 => lut_f_27,
            I1 => lut_f_28,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_30 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_30,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_31 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_31,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_32 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_32,
            I0 => lut_f_30,
            I1 => lut_f_31,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_33 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_33,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_34 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_34,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_35 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_35,
            I0 => lut_f_33,
            I1 => lut_f_34,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_36 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_36,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_37 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_37,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_38 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_38,
            I0 => lut_f_36,
            I1 => lut_f_37,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_39 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_39,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_40 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_40,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_41 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_41,
            I0 => lut_f_39,
            I1 => lut_f_40,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_42 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_42,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_43 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_43,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_44 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_44,
            I0 => lut_f_42,
            I1 => lut_f_43,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_45 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_45,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_46 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_46,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_47 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_47,
            I0 => lut_f_45,
            I1 => lut_f_46,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_48 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_48,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_49 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_49,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_50 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_50,
            I0 => lut_f_48,
            I1 => lut_f_49,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_51 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_51,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_52 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_52,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_53 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_53,
            I0 => lut_f_51,
            I1 => lut_f_52,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_54 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_54,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_55 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_55,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_56 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_56,
            I0 => lut_f_54,
            I1 => lut_f_55,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_57 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_57,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_58 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_58,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_59 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_59,
            I0 => lut_f_57,
            I1 => lut_f_58,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_60 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_60,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_61 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_61,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_62 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_62,
            I0 => lut_f_60,
            I1 => lut_f_61,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_63 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_63,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_64 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_64,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_65 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_65,
            I0 => lut_f_63,
            I1 => lut_f_64,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_66 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_66,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_67 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_67,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_68 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_68,
            I0 => lut_f_66,
            I1 => lut_f_67,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_69 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_69,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_70 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_70,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_71 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_71,
            I0 => lut_f_69,
            I1 => lut_f_70,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_72 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_72,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_73 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_73,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_74 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_74,
            I0 => lut_f_72,
            I1 => lut_f_73,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_75 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_75,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_76 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_76,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_77 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_77,
            I0 => lut_f_75,
            I1 => lut_f_76,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_78 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_78,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_79 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_79,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_80 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_80,
            I0 => lut_f_78,
            I1 => lut_f_79,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_81 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_81,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_82 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_82,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_83 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_83,
            I0 => lut_f_81,
            I1 => lut_f_82,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_84 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_84,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_85 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_85,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_86 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_86,
            I0 => lut_f_84,
            I1 => lut_f_85,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_87 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_87,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_88 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_88,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_89 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_89,
            I0 => lut_f_87,
            I1 => lut_f_88,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_90 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_90,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_91 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_91,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_92 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_92,
            I0 => lut_f_90,
            I1 => lut_f_91,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_93 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_93,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_94 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_94,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad10_inv
        );

    lut_inst_95 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_95,
            I0 => lut_f_93,
            I1 => lut_f_94,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_96 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_96,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_97 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_97,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_98 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_98,
            I0 => lut_f_96,
            I1 => lut_f_97,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_99 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_99,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_100 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_100,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_101 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_101,
            I0 => lut_f_99,
            I1 => lut_f_100,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_102 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_102,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_103 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_103,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_104 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_104,
            I0 => lut_f_102,
            I1 => lut_f_103,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_105 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_105,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_106 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_106,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_107 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_107,
            I0 => lut_f_105,
            I1 => lut_f_106,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_108 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_108,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_109 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_109,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_110 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_110,
            I0 => lut_f_108,
            I1 => lut_f_109,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_111 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_111,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_112 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_112,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_113 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_113,
            I0 => lut_f_111,
            I1 => lut_f_112,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_114 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_114,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_115 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_115,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_116 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_116,
            I0 => lut_f_114,
            I1 => lut_f_115,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_117 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_117,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_118 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_118,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_119 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_119,
            I0 => lut_f_117,
            I1 => lut_f_118,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_120 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_120,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_121 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_121,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_122 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_122,
            I0 => lut_f_120,
            I1 => lut_f_121,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_123 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_123,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_124 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_124,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_125 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_125,
            I0 => lut_f_123,
            I1 => lut_f_124,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_126 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_126,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_127 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_127,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_128 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_128,
            I0 => lut_f_126,
            I1 => lut_f_127,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_129 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_129,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_130 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_130,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_131 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_131,
            I0 => lut_f_129,
            I1 => lut_f_130,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_132 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_132,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_133 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_133,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_134 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_134,
            I0 => lut_f_132,
            I1 => lut_f_133,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_135 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_135,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_136 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_136,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_137 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_137,
            I0 => lut_f_135,
            I1 => lut_f_136,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_138 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_138,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_139 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_139,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_140 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_140,
            I0 => lut_f_138,
            I1 => lut_f_139,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_141 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_141,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_142 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_142,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_143 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_143,
            I0 => lut_f_141,
            I1 => lut_f_142,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_144 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_144,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_145 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_145,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_146 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_146,
            I0 => lut_f_144,
            I1 => lut_f_145,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_147 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_147,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_148 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_148,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_149 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_149,
            I0 => lut_f_147,
            I1 => lut_f_148,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_150 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_150,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_151 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_151,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_152 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_152,
            I0 => lut_f_150,
            I1 => lut_f_151,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_153 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_153,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_154 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_154,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_155 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_155,
            I0 => lut_f_153,
            I1 => lut_f_154,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_156 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_156,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_157 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_157,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_158 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_158,
            I0 => lut_f_156,
            I1 => lut_f_157,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_159 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_159,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_160 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_160,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_161 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_161,
            I0 => lut_f_159,
            I1 => lut_f_160,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_162 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_162,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_163 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_163,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_164 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_164,
            I0 => lut_f_162,
            I1 => lut_f_163,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_165 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_165,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_166 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_166,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_167 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_167,
            I0 => lut_f_165,
            I1 => lut_f_166,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_168 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_168,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_169 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_169,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_170 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_170,
            I0 => lut_f_168,
            I1 => lut_f_169,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_171 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_171,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_172 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_172,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_173 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_173,
            I0 => lut_f_171,
            I1 => lut_f_172,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_174 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_174,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_175 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_175,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_176 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_176,
            I0 => lut_f_174,
            I1 => lut_f_175,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_177 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_177,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_178 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_178,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_179 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_179,
            I0 => lut_f_177,
            I1 => lut_f_178,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_180 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_180,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_181 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_181,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_182 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_182,
            I0 => lut_f_180,
            I1 => lut_f_181,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_183 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_183,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_184 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_184,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_185 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_185,
            I0 => lut_f_183,
            I1 => lut_f_184,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_186 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_186,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_187 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_187,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_188 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_188,
            I0 => lut_f_186,
            I1 => lut_f_187,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_189 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_189,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_190 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_190,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad10_inv
        );

    lut_inst_191 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_191,
            I0 => lut_f_189,
            I1 => lut_f_190,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_192 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_192,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_193 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_193,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_194 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_194,
            I0 => lut_f_192,
            I1 => lut_f_193,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_195 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_195,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_196 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_196,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_197 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_197,
            I0 => lut_f_195,
            I1 => lut_f_196,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_198 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_198,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_199 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_199,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_200 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_200,
            I0 => lut_f_198,
            I1 => lut_f_199,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_201 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_201,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_202 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_202,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_203 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_203,
            I0 => lut_f_201,
            I1 => lut_f_202,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_204 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_204,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_205 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_205,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_206 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_206,
            I0 => lut_f_204,
            I1 => lut_f_205,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_207 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_207,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_208 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_208,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_209 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_209,
            I0 => lut_f_207,
            I1 => lut_f_208,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_210 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_210,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_211 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_211,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_212 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_212,
            I0 => lut_f_210,
            I1 => lut_f_211,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_213 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_213,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_214 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_214,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_215 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_215,
            I0 => lut_f_213,
            I1 => lut_f_214,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_216 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_216,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_217 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_217,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_218 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_218,
            I0 => lut_f_216,
            I1 => lut_f_217,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_219 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_219,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_220 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_220,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_221 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_221,
            I0 => lut_f_219,
            I1 => lut_f_220,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_222 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_222,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_223 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_223,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_224 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_224,
            I0 => lut_f_222,
            I1 => lut_f_223,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_225 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_225,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_226 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_226,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_227 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_227,
            I0 => lut_f_225,
            I1 => lut_f_226,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_228 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_228,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_229 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_229,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_230 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_230,
            I0 => lut_f_228,
            I1 => lut_f_229,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_231 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_231,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_232 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_232,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_233 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_233,
            I0 => lut_f_231,
            I1 => lut_f_232,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_234 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_234,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_235 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_235,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_236 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_236,
            I0 => lut_f_234,
            I1 => lut_f_235,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_237 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_237,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_238 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_238,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_239 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_239,
            I0 => lut_f_237,
            I1 => lut_f_238,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_240 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_240,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_241 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_241,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_242 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_242,
            I0 => lut_f_240,
            I1 => lut_f_241,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_243 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_243,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_244 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_244,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_245 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_245,
            I0 => lut_f_243,
            I1 => lut_f_244,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_246 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_246,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_247 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_247,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_248 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_248,
            I0 => lut_f_246,
            I1 => lut_f_247,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_249 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_249,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_250 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_250,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_251 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_251,
            I0 => lut_f_249,
            I1 => lut_f_250,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_252 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_252,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_253 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_253,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_254 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_254,
            I0 => lut_f_252,
            I1 => lut_f_253,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_255 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_255,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_256 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_256,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_257 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_257,
            I0 => lut_f_255,
            I1 => lut_f_256,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_258 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_258,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_259 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_259,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_260 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_260,
            I0 => lut_f_258,
            I1 => lut_f_259,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_261 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_261,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_262 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_262,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_263 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_263,
            I0 => lut_f_261,
            I1 => lut_f_262,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_264 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_264,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_265 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_265,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_266 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_266,
            I0 => lut_f_264,
            I1 => lut_f_265,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_267 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_267,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_268 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_268,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_269 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_269,
            I0 => lut_f_267,
            I1 => lut_f_268,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_270 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_270,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_271 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_271,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_272 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_272,
            I0 => lut_f_270,
            I1 => lut_f_271,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_273 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_273,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_274 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_274,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_275 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_275,
            I0 => lut_f_273,
            I1 => lut_f_274,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_276 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_276,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_277 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_277,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_278 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_278,
            I0 => lut_f_276,
            I1 => lut_f_277,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_279 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_279,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_280 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_280,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_281 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_281,
            I0 => lut_f_279,
            I1 => lut_f_280,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_282 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_282,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_283 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_283,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_284 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_284,
            I0 => lut_f_282,
            I1 => lut_f_283,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_285 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_285,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_286 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_286,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad9_inv,
            I3 => ad(10)
        );

    lut_inst_287 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_287,
            I0 => lut_f_285,
            I1 => lut_f_286,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_288 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_288,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_289 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_289,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_290 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_290,
            I0 => lut_f_288,
            I1 => lut_f_289,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_291 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_291,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_292 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_292,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_293 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_293,
            I0 => lut_f_291,
            I1 => lut_f_292,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_294 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_294,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_295 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_295,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_296 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_296,
            I0 => lut_f_294,
            I1 => lut_f_295,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_297 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_297,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_298 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_298,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_299 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_299,
            I0 => lut_f_297,
            I1 => lut_f_298,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_300 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_300,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_301 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_301,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_302 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_302,
            I0 => lut_f_300,
            I1 => lut_f_301,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_303 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_303,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_304 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_304,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_305 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_305,
            I0 => lut_f_303,
            I1 => lut_f_304,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_306 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_306,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_307 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_307,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_308 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_308,
            I0 => lut_f_306,
            I1 => lut_f_307,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_309 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_309,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_310 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_310,
            I0 => ad7_inv,
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_311 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_311,
            I0 => lut_f_309,
            I1 => lut_f_310,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_312 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_312,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_313 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_313,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_314 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_314,
            I0 => lut_f_312,
            I1 => lut_f_313,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_315 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_315,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_316 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_316,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_317 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_317,
            I0 => lut_f_315,
            I1 => lut_f_316,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_318 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_318,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_319 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_319,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_320 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_320,
            I0 => lut_f_318,
            I1 => lut_f_319,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_321 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_321,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_322 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_322,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_323 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_323,
            I0 => lut_f_321,
            I1 => lut_f_322,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_324 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_324,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_325 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_325,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_326 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_326,
            I0 => lut_f_324,
            I1 => lut_f_325,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_327 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_327,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_328 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_328,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_329 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_329,
            I0 => lut_f_327,
            I1 => lut_f_328,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_330 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_330,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_331 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_331,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_332 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_332,
            I0 => lut_f_330,
            I1 => lut_f_331,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_333 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_333,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_334 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_334,
            I0 => ad(7),
            I1 => ad8_inv,
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_335 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_335,
            I0 => lut_f_333,
            I1 => lut_f_334,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_336 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_336,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_337 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_337,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_338 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_338,
            I0 => lut_f_336,
            I1 => lut_f_337,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_339 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_339,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_340 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_340,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_341 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_341,
            I0 => lut_f_339,
            I1 => lut_f_340,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_342 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_342,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_343 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_343,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_344 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_344,
            I0 => lut_f_342,
            I1 => lut_f_343,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_345 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_345,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_346 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_346,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_347 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_347,
            I0 => lut_f_345,
            I1 => lut_f_346,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_348 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_348,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_349 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_349,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_350 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_350,
            I0 => lut_f_348,
            I1 => lut_f_349,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_351 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_351,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_352 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_352,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_353 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_353,
            I0 => lut_f_351,
            I1 => lut_f_352,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_354 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_354,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_355 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_355,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_356 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_356,
            I0 => lut_f_354,
            I1 => lut_f_355,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_357 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_357,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_358 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_358,
            I0 => ad7_inv,
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_359 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_359,
            I0 => lut_f_357,
            I1 => lut_f_358,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_360 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_360,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_361 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_361,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_362 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_362,
            I0 => lut_f_360,
            I1 => lut_f_361,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_363 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_363,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_364 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_364,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_365 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_365,
            I0 => lut_f_363,
            I1 => lut_f_364,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_366 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_366,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_367 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_367,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_368 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_368,
            I0 => lut_f_366,
            I1 => lut_f_367,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_369 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_369,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_370 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_370,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_371 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_371,
            I0 => lut_f_369,
            I1 => lut_f_370,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_372 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_372,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_373 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_373,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_374 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_374,
            I0 => lut_f_372,
            I1 => lut_f_373,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_375 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_375,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_376 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_376,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_377 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_377,
            I0 => lut_f_375,
            I1 => lut_f_376,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_378 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_378,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_379 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_379,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_380 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_380,
            I0 => lut_f_378,
            I1 => lut_f_379,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    lut_inst_381 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_381,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_382 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_382,
            I0 => ad(7),
            I1 => ad(8),
            I2 => ad(9),
            I3 => ad(10)
        );

    lut_inst_383 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_383,
            I0 => lut_f_381,
            I1 => lut_f_382,
            I2 => gw_vcc,
            I3 => gw_vcc
        );

    ram16s_inst_0: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_0_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_2,
            CLK => clk
        );

    ram16s_inst_1: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_1_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_2,
            CLK => clk
        );

    ram16s_inst_2: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_2_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_5,
            CLK => clk
        );

    ram16s_inst_3: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_3_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_5,
            CLK => clk
        );

    ram16s_inst_4: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_4_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_8,
            CLK => clk
        );

    ram16s_inst_5: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_5_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_8,
            CLK => clk
        );

    ram16s_inst_6: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_6_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_11,
            CLK => clk
        );

    ram16s_inst_7: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_7_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_11,
            CLK => clk
        );

    ram16s_inst_8: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_8_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_14,
            CLK => clk
        );

    ram16s_inst_9: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_9_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_14,
            CLK => clk
        );

    ram16s_inst_10: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_10_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_17,
            CLK => clk
        );

    ram16s_inst_11: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_11_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_17,
            CLK => clk
        );

    ram16s_inst_12: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_12_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_20,
            CLK => clk
        );

    ram16s_inst_13: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_13_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_20,
            CLK => clk
        );

    ram16s_inst_14: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_14_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_23,
            CLK => clk
        );

    ram16s_inst_15: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_15_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_23,
            CLK => clk
        );

    ram16s_inst_16: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_16_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_26,
            CLK => clk
        );

    ram16s_inst_17: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_17_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_26,
            CLK => clk
        );

    ram16s_inst_18: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_18_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_29,
            CLK => clk
        );

    ram16s_inst_19: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_19_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_29,
            CLK => clk
        );

    ram16s_inst_20: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_20_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_32,
            CLK => clk
        );

    ram16s_inst_21: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_21_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_32,
            CLK => clk
        );

    ram16s_inst_22: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_22_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_35,
            CLK => clk
        );

    ram16s_inst_23: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_23_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_35,
            CLK => clk
        );

    ram16s_inst_24: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_24_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_38,
            CLK => clk
        );

    ram16s_inst_25: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_25_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_38,
            CLK => clk
        );

    ram16s_inst_26: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_26_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_41,
            CLK => clk
        );

    ram16s_inst_27: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_27_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_41,
            CLK => clk
        );

    ram16s_inst_28: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_28_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_44,
            CLK => clk
        );

    ram16s_inst_29: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_29_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_44,
            CLK => clk
        );

    ram16s_inst_30: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_30_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_47,
            CLK => clk
        );

    ram16s_inst_31: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_31_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_47,
            CLK => clk
        );

    ram16s_inst_32: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_32_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_50,
            CLK => clk
        );

    ram16s_inst_33: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_33_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_50,
            CLK => clk
        );

    ram16s_inst_34: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_34_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_53,
            CLK => clk
        );

    ram16s_inst_35: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_35_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_53,
            CLK => clk
        );

    ram16s_inst_36: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_36_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_56,
            CLK => clk
        );

    ram16s_inst_37: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_37_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_56,
            CLK => clk
        );

    ram16s_inst_38: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_38_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_59,
            CLK => clk
        );

    ram16s_inst_39: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_39_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_59,
            CLK => clk
        );

    ram16s_inst_40: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_40_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_62,
            CLK => clk
        );

    ram16s_inst_41: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_41_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_62,
            CLK => clk
        );

    ram16s_inst_42: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_42_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_65,
            CLK => clk
        );

    ram16s_inst_43: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_43_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_65,
            CLK => clk
        );

    ram16s_inst_44: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_44_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_68,
            CLK => clk
        );

    ram16s_inst_45: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_45_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_68,
            CLK => clk
        );

    ram16s_inst_46: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_46_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_71,
            CLK => clk
        );

    ram16s_inst_47: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_47_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_71,
            CLK => clk
        );

    ram16s_inst_48: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_48_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_74,
            CLK => clk
        );

    ram16s_inst_49: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_49_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_74,
            CLK => clk
        );

    ram16s_inst_50: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_50_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_77,
            CLK => clk
        );

    ram16s_inst_51: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_51_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_77,
            CLK => clk
        );

    ram16s_inst_52: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_52_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_80,
            CLK => clk
        );

    ram16s_inst_53: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_53_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_80,
            CLK => clk
        );

    ram16s_inst_54: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_54_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_83,
            CLK => clk
        );

    ram16s_inst_55: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_55_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_83,
            CLK => clk
        );

    ram16s_inst_56: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_56_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_86,
            CLK => clk
        );

    ram16s_inst_57: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_57_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_86,
            CLK => clk
        );

    ram16s_inst_58: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_58_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_89,
            CLK => clk
        );

    ram16s_inst_59: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_59_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_89,
            CLK => clk
        );

    ram16s_inst_60: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_60_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_92,
            CLK => clk
        );

    ram16s_inst_61: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_61_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_92,
            CLK => clk
        );

    ram16s_inst_62: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_62_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_95,
            CLK => clk
        );

    ram16s_inst_63: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_63_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_95,
            CLK => clk
        );

    ram16s_inst_64: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_64_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_98,
            CLK => clk
        );

    ram16s_inst_65: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_65_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_98,
            CLK => clk
        );

    ram16s_inst_66: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_66_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_101,
            CLK => clk
        );

    ram16s_inst_67: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_67_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_101,
            CLK => clk
        );

    ram16s_inst_68: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_68_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_104,
            CLK => clk
        );

    ram16s_inst_69: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_69_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_104,
            CLK => clk
        );

    ram16s_inst_70: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_70_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_107,
            CLK => clk
        );

    ram16s_inst_71: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_71_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_107,
            CLK => clk
        );

    ram16s_inst_72: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_72_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_110,
            CLK => clk
        );

    ram16s_inst_73: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_73_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_110,
            CLK => clk
        );

    ram16s_inst_74: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_74_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_113,
            CLK => clk
        );

    ram16s_inst_75: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_75_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_113,
            CLK => clk
        );

    ram16s_inst_76: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_76_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_116,
            CLK => clk
        );

    ram16s_inst_77: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_77_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_116,
            CLK => clk
        );

    ram16s_inst_78: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_78_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_119,
            CLK => clk
        );

    ram16s_inst_79: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_79_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_119,
            CLK => clk
        );

    ram16s_inst_80: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_80_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_122,
            CLK => clk
        );

    ram16s_inst_81: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_81_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_122,
            CLK => clk
        );

    ram16s_inst_82: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_82_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_125,
            CLK => clk
        );

    ram16s_inst_83: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_83_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_125,
            CLK => clk
        );

    ram16s_inst_84: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_84_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_128,
            CLK => clk
        );

    ram16s_inst_85: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_85_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_128,
            CLK => clk
        );

    ram16s_inst_86: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_86_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_131,
            CLK => clk
        );

    ram16s_inst_87: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_87_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_131,
            CLK => clk
        );

    ram16s_inst_88: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_88_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_134,
            CLK => clk
        );

    ram16s_inst_89: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_89_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_134,
            CLK => clk
        );

    ram16s_inst_90: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_90_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_137,
            CLK => clk
        );

    ram16s_inst_91: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_91_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_137,
            CLK => clk
        );

    ram16s_inst_92: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_92_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_140,
            CLK => clk
        );

    ram16s_inst_93: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_93_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_140,
            CLK => clk
        );

    ram16s_inst_94: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_94_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_143,
            CLK => clk
        );

    ram16s_inst_95: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_95_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_143,
            CLK => clk
        );

    ram16s_inst_96: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_96_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_146,
            CLK => clk
        );

    ram16s_inst_97: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_97_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_146,
            CLK => clk
        );

    ram16s_inst_98: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_98_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_149,
            CLK => clk
        );

    ram16s_inst_99: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_99_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_149,
            CLK => clk
        );

    ram16s_inst_100: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_100_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_152,
            CLK => clk
        );

    ram16s_inst_101: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_101_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_152,
            CLK => clk
        );

    ram16s_inst_102: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_102_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_155,
            CLK => clk
        );

    ram16s_inst_103: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_103_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_155,
            CLK => clk
        );

    ram16s_inst_104: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_104_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_158,
            CLK => clk
        );

    ram16s_inst_105: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_105_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_158,
            CLK => clk
        );

    ram16s_inst_106: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_106_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_161,
            CLK => clk
        );

    ram16s_inst_107: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_107_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_161,
            CLK => clk
        );

    ram16s_inst_108: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_108_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_164,
            CLK => clk
        );

    ram16s_inst_109: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_109_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_164,
            CLK => clk
        );

    ram16s_inst_110: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_110_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_167,
            CLK => clk
        );

    ram16s_inst_111: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_111_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_167,
            CLK => clk
        );

    ram16s_inst_112: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_112_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_170,
            CLK => clk
        );

    ram16s_inst_113: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_113_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_170,
            CLK => clk
        );

    ram16s_inst_114: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_114_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_173,
            CLK => clk
        );

    ram16s_inst_115: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_115_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_173,
            CLK => clk
        );

    ram16s_inst_116: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_116_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_176,
            CLK => clk
        );

    ram16s_inst_117: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_117_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_176,
            CLK => clk
        );

    ram16s_inst_118: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_118_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_179,
            CLK => clk
        );

    ram16s_inst_119: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_119_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_179,
            CLK => clk
        );

    ram16s_inst_120: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_120_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_182,
            CLK => clk
        );

    ram16s_inst_121: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_121_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_182,
            CLK => clk
        );

    ram16s_inst_122: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_122_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_185,
            CLK => clk
        );

    ram16s_inst_123: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_123_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_185,
            CLK => clk
        );

    ram16s_inst_124: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_124_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_188,
            CLK => clk
        );

    ram16s_inst_125: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_125_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_188,
            CLK => clk
        );

    ram16s_inst_126: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_126_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_191,
            CLK => clk
        );

    ram16s_inst_127: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_127_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_191,
            CLK => clk
        );

    ram16s_inst_128: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_128_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_194,
            CLK => clk
        );

    ram16s_inst_129: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_129_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_194,
            CLK => clk
        );

    ram16s_inst_130: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_130_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_197,
            CLK => clk
        );

    ram16s_inst_131: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_131_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_197,
            CLK => clk
        );

    ram16s_inst_132: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_132_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_200,
            CLK => clk
        );

    ram16s_inst_133: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_133_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_200,
            CLK => clk
        );

    ram16s_inst_134: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_134_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_203,
            CLK => clk
        );

    ram16s_inst_135: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_135_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_203,
            CLK => clk
        );

    ram16s_inst_136: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_136_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_206,
            CLK => clk
        );

    ram16s_inst_137: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_137_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_206,
            CLK => clk
        );

    ram16s_inst_138: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_138_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_209,
            CLK => clk
        );

    ram16s_inst_139: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_139_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_209,
            CLK => clk
        );

    ram16s_inst_140: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_140_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_212,
            CLK => clk
        );

    ram16s_inst_141: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_141_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_212,
            CLK => clk
        );

    ram16s_inst_142: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_142_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_215,
            CLK => clk
        );

    ram16s_inst_143: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_143_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_215,
            CLK => clk
        );

    ram16s_inst_144: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_144_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_218,
            CLK => clk
        );

    ram16s_inst_145: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_145_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_218,
            CLK => clk
        );

    ram16s_inst_146: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_146_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_221,
            CLK => clk
        );

    ram16s_inst_147: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_147_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_221,
            CLK => clk
        );

    ram16s_inst_148: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_148_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_224,
            CLK => clk
        );

    ram16s_inst_149: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_149_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_224,
            CLK => clk
        );

    ram16s_inst_150: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_150_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_227,
            CLK => clk
        );

    ram16s_inst_151: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_151_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_227,
            CLK => clk
        );

    ram16s_inst_152: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_152_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_230,
            CLK => clk
        );

    ram16s_inst_153: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_153_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_230,
            CLK => clk
        );

    ram16s_inst_154: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_154_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_233,
            CLK => clk
        );

    ram16s_inst_155: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_155_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_233,
            CLK => clk
        );

    ram16s_inst_156: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_156_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_236,
            CLK => clk
        );

    ram16s_inst_157: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_157_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_236,
            CLK => clk
        );

    ram16s_inst_158: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_158_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_239,
            CLK => clk
        );

    ram16s_inst_159: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_159_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_239,
            CLK => clk
        );

    ram16s_inst_160: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_160_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_242,
            CLK => clk
        );

    ram16s_inst_161: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_161_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_242,
            CLK => clk
        );

    ram16s_inst_162: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_162_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_245,
            CLK => clk
        );

    ram16s_inst_163: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_163_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_245,
            CLK => clk
        );

    ram16s_inst_164: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_164_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_248,
            CLK => clk
        );

    ram16s_inst_165: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_165_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_248,
            CLK => clk
        );

    ram16s_inst_166: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_166_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_251,
            CLK => clk
        );

    ram16s_inst_167: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_167_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_251,
            CLK => clk
        );

    ram16s_inst_168: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_168_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_254,
            CLK => clk
        );

    ram16s_inst_169: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_169_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_254,
            CLK => clk
        );

    ram16s_inst_170: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_170_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_257,
            CLK => clk
        );

    ram16s_inst_171: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_171_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_257,
            CLK => clk
        );

    ram16s_inst_172: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_172_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_260,
            CLK => clk
        );

    ram16s_inst_173: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_173_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_260,
            CLK => clk
        );

    ram16s_inst_174: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_174_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_263,
            CLK => clk
        );

    ram16s_inst_175: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_175_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_263,
            CLK => clk
        );

    ram16s_inst_176: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_176_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_266,
            CLK => clk
        );

    ram16s_inst_177: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_177_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_266,
            CLK => clk
        );

    ram16s_inst_178: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_178_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_269,
            CLK => clk
        );

    ram16s_inst_179: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_179_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_269,
            CLK => clk
        );

    ram16s_inst_180: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_180_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_272,
            CLK => clk
        );

    ram16s_inst_181: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_181_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_272,
            CLK => clk
        );

    ram16s_inst_182: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_182_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_275,
            CLK => clk
        );

    ram16s_inst_183: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_183_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_275,
            CLK => clk
        );

    ram16s_inst_184: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_184_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_278,
            CLK => clk
        );

    ram16s_inst_185: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_185_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_278,
            CLK => clk
        );

    ram16s_inst_186: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_186_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_281,
            CLK => clk
        );

    ram16s_inst_187: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_187_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_281,
            CLK => clk
        );

    ram16s_inst_188: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_188_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_284,
            CLK => clk
        );

    ram16s_inst_189: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_189_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_284,
            CLK => clk
        );

    ram16s_inst_190: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_190_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_287,
            CLK => clk
        );

    ram16s_inst_191: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_191_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_287,
            CLK => clk
        );

    ram16s_inst_192: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_192_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_290,
            CLK => clk
        );

    ram16s_inst_193: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_193_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_290,
            CLK => clk
        );

    ram16s_inst_194: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_194_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_293,
            CLK => clk
        );

    ram16s_inst_195: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_195_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_293,
            CLK => clk
        );

    ram16s_inst_196: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_196_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_296,
            CLK => clk
        );

    ram16s_inst_197: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_197_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_296,
            CLK => clk
        );

    ram16s_inst_198: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_198_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_299,
            CLK => clk
        );

    ram16s_inst_199: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_199_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_299,
            CLK => clk
        );

    ram16s_inst_200: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_200_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_302,
            CLK => clk
        );

    ram16s_inst_201: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_201_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_302,
            CLK => clk
        );

    ram16s_inst_202: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_202_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_305,
            CLK => clk
        );

    ram16s_inst_203: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_203_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_305,
            CLK => clk
        );

    ram16s_inst_204: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_204_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_308,
            CLK => clk
        );

    ram16s_inst_205: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_205_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_308,
            CLK => clk
        );

    ram16s_inst_206: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_206_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_311,
            CLK => clk
        );

    ram16s_inst_207: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_207_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_311,
            CLK => clk
        );

    ram16s_inst_208: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_208_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_314,
            CLK => clk
        );

    ram16s_inst_209: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_209_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_314,
            CLK => clk
        );

    ram16s_inst_210: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_210_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_317,
            CLK => clk
        );

    ram16s_inst_211: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_211_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_317,
            CLK => clk
        );

    ram16s_inst_212: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_212_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_320,
            CLK => clk
        );

    ram16s_inst_213: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_213_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_320,
            CLK => clk
        );

    ram16s_inst_214: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_214_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_323,
            CLK => clk
        );

    ram16s_inst_215: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_215_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_323,
            CLK => clk
        );

    ram16s_inst_216: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_216_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_326,
            CLK => clk
        );

    ram16s_inst_217: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_217_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_326,
            CLK => clk
        );

    ram16s_inst_218: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_218_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_329,
            CLK => clk
        );

    ram16s_inst_219: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_219_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_329,
            CLK => clk
        );

    ram16s_inst_220: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_220_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_332,
            CLK => clk
        );

    ram16s_inst_221: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_221_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_332,
            CLK => clk
        );

    ram16s_inst_222: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_222_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_335,
            CLK => clk
        );

    ram16s_inst_223: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_223_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_335,
            CLK => clk
        );

    ram16s_inst_224: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_224_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_338,
            CLK => clk
        );

    ram16s_inst_225: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_225_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_338,
            CLK => clk
        );

    ram16s_inst_226: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_226_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_341,
            CLK => clk
        );

    ram16s_inst_227: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_227_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_341,
            CLK => clk
        );

    ram16s_inst_228: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_228_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_344,
            CLK => clk
        );

    ram16s_inst_229: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_229_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_344,
            CLK => clk
        );

    ram16s_inst_230: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_230_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_347,
            CLK => clk
        );

    ram16s_inst_231: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_231_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_347,
            CLK => clk
        );

    ram16s_inst_232: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_232_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_350,
            CLK => clk
        );

    ram16s_inst_233: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_233_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_350,
            CLK => clk
        );

    ram16s_inst_234: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_234_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_353,
            CLK => clk
        );

    ram16s_inst_235: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_235_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_353,
            CLK => clk
        );

    ram16s_inst_236: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_236_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_356,
            CLK => clk
        );

    ram16s_inst_237: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_237_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_356,
            CLK => clk
        );

    ram16s_inst_238: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_238_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_359,
            CLK => clk
        );

    ram16s_inst_239: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_239_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_359,
            CLK => clk
        );

    ram16s_inst_240: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_240_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_362,
            CLK => clk
        );

    ram16s_inst_241: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_241_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_362,
            CLK => clk
        );

    ram16s_inst_242: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_242_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_365,
            CLK => clk
        );

    ram16s_inst_243: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_243_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_365,
            CLK => clk
        );

    ram16s_inst_244: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_244_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_368,
            CLK => clk
        );

    ram16s_inst_245: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_245_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_368,
            CLK => clk
        );

    ram16s_inst_246: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_246_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_371,
            CLK => clk
        );

    ram16s_inst_247: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_247_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_371,
            CLK => clk
        );

    ram16s_inst_248: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_248_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_374,
            CLK => clk
        );

    ram16s_inst_249: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_249_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_374,
            CLK => clk
        );

    ram16s_inst_250: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_250_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_377,
            CLK => clk
        );

    ram16s_inst_251: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_251_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_377,
            CLK => clk
        );

    ram16s_inst_252: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_252_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_380,
            CLK => clk
        );

    ram16s_inst_253: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_253_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_380,
            CLK => clk
        );

    ram16s_inst_254: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_254_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_383,
            CLK => clk
        );

    ram16s_inst_255: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_255_dout(7 downto 4),
            DI => di(7 downto 4),
            AD => ad(3 downto 0),
            WRE => lut_f_383,
            CLK => clk
        );

    mux_inst_0: MUX2
        port map (
            O => mux_o_0,
            I0 => ram16s_inst_0_dout(0),
            I1 => ram16s_inst_2_dout(0),
            S0 => ad(4)
        );

    mux_inst_1: MUX2
        port map (
            O => mux_o_1,
            I0 => ram16s_inst_4_dout(0),
            I1 => ram16s_inst_6_dout(0),
            S0 => ad(4)
        );

    mux_inst_2: MUX2
        port map (
            O => mux_o_2,
            I0 => ram16s_inst_8_dout(0),
            I1 => ram16s_inst_10_dout(0),
            S0 => ad(4)
        );

    mux_inst_3: MUX2
        port map (
            O => mux_o_3,
            I0 => ram16s_inst_12_dout(0),
            I1 => ram16s_inst_14_dout(0),
            S0 => ad(4)
        );

    mux_inst_4: MUX2
        port map (
            O => mux_o_4,
            I0 => ram16s_inst_16_dout(0),
            I1 => ram16s_inst_18_dout(0),
            S0 => ad(4)
        );

    mux_inst_5: MUX2
        port map (
            O => mux_o_5,
            I0 => ram16s_inst_20_dout(0),
            I1 => ram16s_inst_22_dout(0),
            S0 => ad(4)
        );

    mux_inst_6: MUX2
        port map (
            O => mux_o_6,
            I0 => ram16s_inst_24_dout(0),
            I1 => ram16s_inst_26_dout(0),
            S0 => ad(4)
        );

    mux_inst_7: MUX2
        port map (
            O => mux_o_7,
            I0 => ram16s_inst_28_dout(0),
            I1 => ram16s_inst_30_dout(0),
            S0 => ad(4)
        );

    mux_inst_8: MUX2
        port map (
            O => mux_o_8,
            I0 => ram16s_inst_32_dout(0),
            I1 => ram16s_inst_34_dout(0),
            S0 => ad(4)
        );

    mux_inst_9: MUX2
        port map (
            O => mux_o_9,
            I0 => ram16s_inst_36_dout(0),
            I1 => ram16s_inst_38_dout(0),
            S0 => ad(4)
        );

    mux_inst_10: MUX2
        port map (
            O => mux_o_10,
            I0 => ram16s_inst_40_dout(0),
            I1 => ram16s_inst_42_dout(0),
            S0 => ad(4)
        );

    mux_inst_11: MUX2
        port map (
            O => mux_o_11,
            I0 => ram16s_inst_44_dout(0),
            I1 => ram16s_inst_46_dout(0),
            S0 => ad(4)
        );

    mux_inst_12: MUX2
        port map (
            O => mux_o_12,
            I0 => ram16s_inst_48_dout(0),
            I1 => ram16s_inst_50_dout(0),
            S0 => ad(4)
        );

    mux_inst_13: MUX2
        port map (
            O => mux_o_13,
            I0 => ram16s_inst_52_dout(0),
            I1 => ram16s_inst_54_dout(0),
            S0 => ad(4)
        );

    mux_inst_14: MUX2
        port map (
            O => mux_o_14,
            I0 => ram16s_inst_56_dout(0),
            I1 => ram16s_inst_58_dout(0),
            S0 => ad(4)
        );

    mux_inst_15: MUX2
        port map (
            O => mux_o_15,
            I0 => ram16s_inst_60_dout(0),
            I1 => ram16s_inst_62_dout(0),
            S0 => ad(4)
        );

    mux_inst_16: MUX2
        port map (
            O => mux_o_16,
            I0 => ram16s_inst_64_dout(0),
            I1 => ram16s_inst_66_dout(0),
            S0 => ad(4)
        );

    mux_inst_17: MUX2
        port map (
            O => mux_o_17,
            I0 => ram16s_inst_68_dout(0),
            I1 => ram16s_inst_70_dout(0),
            S0 => ad(4)
        );

    mux_inst_18: MUX2
        port map (
            O => mux_o_18,
            I0 => ram16s_inst_72_dout(0),
            I1 => ram16s_inst_74_dout(0),
            S0 => ad(4)
        );

    mux_inst_19: MUX2
        port map (
            O => mux_o_19,
            I0 => ram16s_inst_76_dout(0),
            I1 => ram16s_inst_78_dout(0),
            S0 => ad(4)
        );

    mux_inst_20: MUX2
        port map (
            O => mux_o_20,
            I0 => ram16s_inst_80_dout(0),
            I1 => ram16s_inst_82_dout(0),
            S0 => ad(4)
        );

    mux_inst_21: MUX2
        port map (
            O => mux_o_21,
            I0 => ram16s_inst_84_dout(0),
            I1 => ram16s_inst_86_dout(0),
            S0 => ad(4)
        );

    mux_inst_22: MUX2
        port map (
            O => mux_o_22,
            I0 => ram16s_inst_88_dout(0),
            I1 => ram16s_inst_90_dout(0),
            S0 => ad(4)
        );

    mux_inst_23: MUX2
        port map (
            O => mux_o_23,
            I0 => ram16s_inst_92_dout(0),
            I1 => ram16s_inst_94_dout(0),
            S0 => ad(4)
        );

    mux_inst_24: MUX2
        port map (
            O => mux_o_24,
            I0 => ram16s_inst_96_dout(0),
            I1 => ram16s_inst_98_dout(0),
            S0 => ad(4)
        );

    mux_inst_25: MUX2
        port map (
            O => mux_o_25,
            I0 => ram16s_inst_100_dout(0),
            I1 => ram16s_inst_102_dout(0),
            S0 => ad(4)
        );

    mux_inst_26: MUX2
        port map (
            O => mux_o_26,
            I0 => ram16s_inst_104_dout(0),
            I1 => ram16s_inst_106_dout(0),
            S0 => ad(4)
        );

    mux_inst_27: MUX2
        port map (
            O => mux_o_27,
            I0 => ram16s_inst_108_dout(0),
            I1 => ram16s_inst_110_dout(0),
            S0 => ad(4)
        );

    mux_inst_28: MUX2
        port map (
            O => mux_o_28,
            I0 => ram16s_inst_112_dout(0),
            I1 => ram16s_inst_114_dout(0),
            S0 => ad(4)
        );

    mux_inst_29: MUX2
        port map (
            O => mux_o_29,
            I0 => ram16s_inst_116_dout(0),
            I1 => ram16s_inst_118_dout(0),
            S0 => ad(4)
        );

    mux_inst_30: MUX2
        port map (
            O => mux_o_30,
            I0 => ram16s_inst_120_dout(0),
            I1 => ram16s_inst_122_dout(0),
            S0 => ad(4)
        );

    mux_inst_31: MUX2
        port map (
            O => mux_o_31,
            I0 => ram16s_inst_124_dout(0),
            I1 => ram16s_inst_126_dout(0),
            S0 => ad(4)
        );

    mux_inst_32: MUX2
        port map (
            O => mux_o_32,
            I0 => ram16s_inst_128_dout(0),
            I1 => ram16s_inst_130_dout(0),
            S0 => ad(4)
        );

    mux_inst_33: MUX2
        port map (
            O => mux_o_33,
            I0 => ram16s_inst_132_dout(0),
            I1 => ram16s_inst_134_dout(0),
            S0 => ad(4)
        );

    mux_inst_34: MUX2
        port map (
            O => mux_o_34,
            I0 => ram16s_inst_136_dout(0),
            I1 => ram16s_inst_138_dout(0),
            S0 => ad(4)
        );

    mux_inst_35: MUX2
        port map (
            O => mux_o_35,
            I0 => ram16s_inst_140_dout(0),
            I1 => ram16s_inst_142_dout(0),
            S0 => ad(4)
        );

    mux_inst_36: MUX2
        port map (
            O => mux_o_36,
            I0 => ram16s_inst_144_dout(0),
            I1 => ram16s_inst_146_dout(0),
            S0 => ad(4)
        );

    mux_inst_37: MUX2
        port map (
            O => mux_o_37,
            I0 => ram16s_inst_148_dout(0),
            I1 => ram16s_inst_150_dout(0),
            S0 => ad(4)
        );

    mux_inst_38: MUX2
        port map (
            O => mux_o_38,
            I0 => ram16s_inst_152_dout(0),
            I1 => ram16s_inst_154_dout(0),
            S0 => ad(4)
        );

    mux_inst_39: MUX2
        port map (
            O => mux_o_39,
            I0 => ram16s_inst_156_dout(0),
            I1 => ram16s_inst_158_dout(0),
            S0 => ad(4)
        );

    mux_inst_40: MUX2
        port map (
            O => mux_o_40,
            I0 => ram16s_inst_160_dout(0),
            I1 => ram16s_inst_162_dout(0),
            S0 => ad(4)
        );

    mux_inst_41: MUX2
        port map (
            O => mux_o_41,
            I0 => ram16s_inst_164_dout(0),
            I1 => ram16s_inst_166_dout(0),
            S0 => ad(4)
        );

    mux_inst_42: MUX2
        port map (
            O => mux_o_42,
            I0 => ram16s_inst_168_dout(0),
            I1 => ram16s_inst_170_dout(0),
            S0 => ad(4)
        );

    mux_inst_43: MUX2
        port map (
            O => mux_o_43,
            I0 => ram16s_inst_172_dout(0),
            I1 => ram16s_inst_174_dout(0),
            S0 => ad(4)
        );

    mux_inst_44: MUX2
        port map (
            O => mux_o_44,
            I0 => ram16s_inst_176_dout(0),
            I1 => ram16s_inst_178_dout(0),
            S0 => ad(4)
        );

    mux_inst_45: MUX2
        port map (
            O => mux_o_45,
            I0 => ram16s_inst_180_dout(0),
            I1 => ram16s_inst_182_dout(0),
            S0 => ad(4)
        );

    mux_inst_46: MUX2
        port map (
            O => mux_o_46,
            I0 => ram16s_inst_184_dout(0),
            I1 => ram16s_inst_186_dout(0),
            S0 => ad(4)
        );

    mux_inst_47: MUX2
        port map (
            O => mux_o_47,
            I0 => ram16s_inst_188_dout(0),
            I1 => ram16s_inst_190_dout(0),
            S0 => ad(4)
        );

    mux_inst_48: MUX2
        port map (
            O => mux_o_48,
            I0 => ram16s_inst_192_dout(0),
            I1 => ram16s_inst_194_dout(0),
            S0 => ad(4)
        );

    mux_inst_49: MUX2
        port map (
            O => mux_o_49,
            I0 => ram16s_inst_196_dout(0),
            I1 => ram16s_inst_198_dout(0),
            S0 => ad(4)
        );

    mux_inst_50: MUX2
        port map (
            O => mux_o_50,
            I0 => ram16s_inst_200_dout(0),
            I1 => ram16s_inst_202_dout(0),
            S0 => ad(4)
        );

    mux_inst_51: MUX2
        port map (
            O => mux_o_51,
            I0 => ram16s_inst_204_dout(0),
            I1 => ram16s_inst_206_dout(0),
            S0 => ad(4)
        );

    mux_inst_52: MUX2
        port map (
            O => mux_o_52,
            I0 => ram16s_inst_208_dout(0),
            I1 => ram16s_inst_210_dout(0),
            S0 => ad(4)
        );

    mux_inst_53: MUX2
        port map (
            O => mux_o_53,
            I0 => ram16s_inst_212_dout(0),
            I1 => ram16s_inst_214_dout(0),
            S0 => ad(4)
        );

    mux_inst_54: MUX2
        port map (
            O => mux_o_54,
            I0 => ram16s_inst_216_dout(0),
            I1 => ram16s_inst_218_dout(0),
            S0 => ad(4)
        );

    mux_inst_55: MUX2
        port map (
            O => mux_o_55,
            I0 => ram16s_inst_220_dout(0),
            I1 => ram16s_inst_222_dout(0),
            S0 => ad(4)
        );

    mux_inst_56: MUX2
        port map (
            O => mux_o_56,
            I0 => ram16s_inst_224_dout(0),
            I1 => ram16s_inst_226_dout(0),
            S0 => ad(4)
        );

    mux_inst_57: MUX2
        port map (
            O => mux_o_57,
            I0 => ram16s_inst_228_dout(0),
            I1 => ram16s_inst_230_dout(0),
            S0 => ad(4)
        );

    mux_inst_58: MUX2
        port map (
            O => mux_o_58,
            I0 => ram16s_inst_232_dout(0),
            I1 => ram16s_inst_234_dout(0),
            S0 => ad(4)
        );

    mux_inst_59: MUX2
        port map (
            O => mux_o_59,
            I0 => ram16s_inst_236_dout(0),
            I1 => ram16s_inst_238_dout(0),
            S0 => ad(4)
        );

    mux_inst_60: MUX2
        port map (
            O => mux_o_60,
            I0 => ram16s_inst_240_dout(0),
            I1 => ram16s_inst_242_dout(0),
            S0 => ad(4)
        );

    mux_inst_61: MUX2
        port map (
            O => mux_o_61,
            I0 => ram16s_inst_244_dout(0),
            I1 => ram16s_inst_246_dout(0),
            S0 => ad(4)
        );

    mux_inst_62: MUX2
        port map (
            O => mux_o_62,
            I0 => ram16s_inst_248_dout(0),
            I1 => ram16s_inst_250_dout(0),
            S0 => ad(4)
        );

    mux_inst_63: MUX2
        port map (
            O => mux_o_63,
            I0 => ram16s_inst_252_dout(0),
            I1 => ram16s_inst_254_dout(0),
            S0 => ad(4)
        );

    mux_inst_64: MUX2
        port map (
            O => mux_o_64,
            I0 => mux_o_0,
            I1 => mux_o_1,
            S0 => ad(5)
        );

    mux_inst_65: MUX2
        port map (
            O => mux_o_65,
            I0 => mux_o_2,
            I1 => mux_o_3,
            S0 => ad(5)
        );

    mux_inst_66: MUX2
        port map (
            O => mux_o_66,
            I0 => mux_o_4,
            I1 => mux_o_5,
            S0 => ad(5)
        );

    mux_inst_67: MUX2
        port map (
            O => mux_o_67,
            I0 => mux_o_6,
            I1 => mux_o_7,
            S0 => ad(5)
        );

    mux_inst_68: MUX2
        port map (
            O => mux_o_68,
            I0 => mux_o_8,
            I1 => mux_o_9,
            S0 => ad(5)
        );

    mux_inst_69: MUX2
        port map (
            O => mux_o_69,
            I0 => mux_o_10,
            I1 => mux_o_11,
            S0 => ad(5)
        );

    mux_inst_70: MUX2
        port map (
            O => mux_o_70,
            I0 => mux_o_12,
            I1 => mux_o_13,
            S0 => ad(5)
        );

    mux_inst_71: MUX2
        port map (
            O => mux_o_71,
            I0 => mux_o_14,
            I1 => mux_o_15,
            S0 => ad(5)
        );

    mux_inst_72: MUX2
        port map (
            O => mux_o_72,
            I0 => mux_o_16,
            I1 => mux_o_17,
            S0 => ad(5)
        );

    mux_inst_73: MUX2
        port map (
            O => mux_o_73,
            I0 => mux_o_18,
            I1 => mux_o_19,
            S0 => ad(5)
        );

    mux_inst_74: MUX2
        port map (
            O => mux_o_74,
            I0 => mux_o_20,
            I1 => mux_o_21,
            S0 => ad(5)
        );

    mux_inst_75: MUX2
        port map (
            O => mux_o_75,
            I0 => mux_o_22,
            I1 => mux_o_23,
            S0 => ad(5)
        );

    mux_inst_76: MUX2
        port map (
            O => mux_o_76,
            I0 => mux_o_24,
            I1 => mux_o_25,
            S0 => ad(5)
        );

    mux_inst_77: MUX2
        port map (
            O => mux_o_77,
            I0 => mux_o_26,
            I1 => mux_o_27,
            S0 => ad(5)
        );

    mux_inst_78: MUX2
        port map (
            O => mux_o_78,
            I0 => mux_o_28,
            I1 => mux_o_29,
            S0 => ad(5)
        );

    mux_inst_79: MUX2
        port map (
            O => mux_o_79,
            I0 => mux_o_30,
            I1 => mux_o_31,
            S0 => ad(5)
        );

    mux_inst_80: MUX2
        port map (
            O => mux_o_80,
            I0 => mux_o_32,
            I1 => mux_o_33,
            S0 => ad(5)
        );

    mux_inst_81: MUX2
        port map (
            O => mux_o_81,
            I0 => mux_o_34,
            I1 => mux_o_35,
            S0 => ad(5)
        );

    mux_inst_82: MUX2
        port map (
            O => mux_o_82,
            I0 => mux_o_36,
            I1 => mux_o_37,
            S0 => ad(5)
        );

    mux_inst_83: MUX2
        port map (
            O => mux_o_83,
            I0 => mux_o_38,
            I1 => mux_o_39,
            S0 => ad(5)
        );

    mux_inst_84: MUX2
        port map (
            O => mux_o_84,
            I0 => mux_o_40,
            I1 => mux_o_41,
            S0 => ad(5)
        );

    mux_inst_85: MUX2
        port map (
            O => mux_o_85,
            I0 => mux_o_42,
            I1 => mux_o_43,
            S0 => ad(5)
        );

    mux_inst_86: MUX2
        port map (
            O => mux_o_86,
            I0 => mux_o_44,
            I1 => mux_o_45,
            S0 => ad(5)
        );

    mux_inst_87: MUX2
        port map (
            O => mux_o_87,
            I0 => mux_o_46,
            I1 => mux_o_47,
            S0 => ad(5)
        );

    mux_inst_88: MUX2
        port map (
            O => mux_o_88,
            I0 => mux_o_48,
            I1 => mux_o_49,
            S0 => ad(5)
        );

    mux_inst_89: MUX2
        port map (
            O => mux_o_89,
            I0 => mux_o_50,
            I1 => mux_o_51,
            S0 => ad(5)
        );

    mux_inst_90: MUX2
        port map (
            O => mux_o_90,
            I0 => mux_o_52,
            I1 => mux_o_53,
            S0 => ad(5)
        );

    mux_inst_91: MUX2
        port map (
            O => mux_o_91,
            I0 => mux_o_54,
            I1 => mux_o_55,
            S0 => ad(5)
        );

    mux_inst_92: MUX2
        port map (
            O => mux_o_92,
            I0 => mux_o_56,
            I1 => mux_o_57,
            S0 => ad(5)
        );

    mux_inst_93: MUX2
        port map (
            O => mux_o_93,
            I0 => mux_o_58,
            I1 => mux_o_59,
            S0 => ad(5)
        );

    mux_inst_94: MUX2
        port map (
            O => mux_o_94,
            I0 => mux_o_60,
            I1 => mux_o_61,
            S0 => ad(5)
        );

    mux_inst_95: MUX2
        port map (
            O => mux_o_95,
            I0 => mux_o_62,
            I1 => mux_o_63,
            S0 => ad(5)
        );

    mux_inst_96: MUX2
        port map (
            O => mux_o_96,
            I0 => mux_o_64,
            I1 => mux_o_65,
            S0 => ad(6)
        );

    mux_inst_97: MUX2
        port map (
            O => mux_o_97,
            I0 => mux_o_66,
            I1 => mux_o_67,
            S0 => ad(6)
        );

    mux_inst_98: MUX2
        port map (
            O => mux_o_98,
            I0 => mux_o_68,
            I1 => mux_o_69,
            S0 => ad(6)
        );

    mux_inst_99: MUX2
        port map (
            O => mux_o_99,
            I0 => mux_o_70,
            I1 => mux_o_71,
            S0 => ad(6)
        );

    mux_inst_100: MUX2
        port map (
            O => mux_o_100,
            I0 => mux_o_72,
            I1 => mux_o_73,
            S0 => ad(6)
        );

    mux_inst_101: MUX2
        port map (
            O => mux_o_101,
            I0 => mux_o_74,
            I1 => mux_o_75,
            S0 => ad(6)
        );

    mux_inst_102: MUX2
        port map (
            O => mux_o_102,
            I0 => mux_o_76,
            I1 => mux_o_77,
            S0 => ad(6)
        );

    mux_inst_103: MUX2
        port map (
            O => mux_o_103,
            I0 => mux_o_78,
            I1 => mux_o_79,
            S0 => ad(6)
        );

    mux_inst_104: MUX2
        port map (
            O => mux_o_104,
            I0 => mux_o_80,
            I1 => mux_o_81,
            S0 => ad(6)
        );

    mux_inst_105: MUX2
        port map (
            O => mux_o_105,
            I0 => mux_o_82,
            I1 => mux_o_83,
            S0 => ad(6)
        );

    mux_inst_106: MUX2
        port map (
            O => mux_o_106,
            I0 => mux_o_84,
            I1 => mux_o_85,
            S0 => ad(6)
        );

    mux_inst_107: MUX2
        port map (
            O => mux_o_107,
            I0 => mux_o_86,
            I1 => mux_o_87,
            S0 => ad(6)
        );

    mux_inst_108: MUX2
        port map (
            O => mux_o_108,
            I0 => mux_o_88,
            I1 => mux_o_89,
            S0 => ad(6)
        );

    mux_inst_109: MUX2
        port map (
            O => mux_o_109,
            I0 => mux_o_90,
            I1 => mux_o_91,
            S0 => ad(6)
        );

    mux_inst_110: MUX2
        port map (
            O => mux_o_110,
            I0 => mux_o_92,
            I1 => mux_o_93,
            S0 => ad(6)
        );

    mux_inst_111: MUX2
        port map (
            O => mux_o_111,
            I0 => mux_o_94,
            I1 => mux_o_95,
            S0 => ad(6)
        );

    mux_inst_112: MUX2
        port map (
            O => mux_o_112,
            I0 => mux_o_96,
            I1 => mux_o_97,
            S0 => ad(7)
        );

    mux_inst_113: MUX2
        port map (
            O => mux_o_113,
            I0 => mux_o_98,
            I1 => mux_o_99,
            S0 => ad(7)
        );

    mux_inst_114: MUX2
        port map (
            O => mux_o_114,
            I0 => mux_o_100,
            I1 => mux_o_101,
            S0 => ad(7)
        );

    mux_inst_115: MUX2
        port map (
            O => mux_o_115,
            I0 => mux_o_102,
            I1 => mux_o_103,
            S0 => ad(7)
        );

    mux_inst_116: MUX2
        port map (
            O => mux_o_116,
            I0 => mux_o_104,
            I1 => mux_o_105,
            S0 => ad(7)
        );

    mux_inst_117: MUX2
        port map (
            O => mux_o_117,
            I0 => mux_o_106,
            I1 => mux_o_107,
            S0 => ad(7)
        );

    mux_inst_118: MUX2
        port map (
            O => mux_o_118,
            I0 => mux_o_108,
            I1 => mux_o_109,
            S0 => ad(7)
        );

    mux_inst_119: MUX2
        port map (
            O => mux_o_119,
            I0 => mux_o_110,
            I1 => mux_o_111,
            S0 => ad(7)
        );

    mux_inst_120: MUX2
        port map (
            O => mux_o_120,
            I0 => mux_o_112,
            I1 => mux_o_113,
            S0 => ad(8)
        );

    mux_inst_121: MUX2
        port map (
            O => mux_o_121,
            I0 => mux_o_114,
            I1 => mux_o_115,
            S0 => ad(8)
        );

    mux_inst_122: MUX2
        port map (
            O => mux_o_122,
            I0 => mux_o_116,
            I1 => mux_o_117,
            S0 => ad(8)
        );

    mux_inst_123: MUX2
        port map (
            O => mux_o_123,
            I0 => mux_o_118,
            I1 => mux_o_119,
            S0 => ad(8)
        );

    mux_inst_124: MUX2
        port map (
            O => mux_o_124,
            I0 => mux_o_120,
            I1 => mux_o_121,
            S0 => ad(9)
        );

    mux_inst_125: MUX2
        port map (
            O => mux_o_125,
            I0 => mux_o_122,
            I1 => mux_o_123,
            S0 => ad(9)
        );

    mux_inst_126: MUX2
        port map (
            O => dout(0),
            I0 => mux_o_124,
            I1 => mux_o_125,
            S0 => ad(10)
        );

    mux_inst_127: MUX2
        port map (
            O => mux_o_127,
            I0 => ram16s_inst_0_dout(1),
            I1 => ram16s_inst_2_dout(1),
            S0 => ad(4)
        );

    mux_inst_128: MUX2
        port map (
            O => mux_o_128,
            I0 => ram16s_inst_4_dout(1),
            I1 => ram16s_inst_6_dout(1),
            S0 => ad(4)
        );

    mux_inst_129: MUX2
        port map (
            O => mux_o_129,
            I0 => ram16s_inst_8_dout(1),
            I1 => ram16s_inst_10_dout(1),
            S0 => ad(4)
        );

    mux_inst_130: MUX2
        port map (
            O => mux_o_130,
            I0 => ram16s_inst_12_dout(1),
            I1 => ram16s_inst_14_dout(1),
            S0 => ad(4)
        );

    mux_inst_131: MUX2
        port map (
            O => mux_o_131,
            I0 => ram16s_inst_16_dout(1),
            I1 => ram16s_inst_18_dout(1),
            S0 => ad(4)
        );

    mux_inst_132: MUX2
        port map (
            O => mux_o_132,
            I0 => ram16s_inst_20_dout(1),
            I1 => ram16s_inst_22_dout(1),
            S0 => ad(4)
        );

    mux_inst_133: MUX2
        port map (
            O => mux_o_133,
            I0 => ram16s_inst_24_dout(1),
            I1 => ram16s_inst_26_dout(1),
            S0 => ad(4)
        );

    mux_inst_134: MUX2
        port map (
            O => mux_o_134,
            I0 => ram16s_inst_28_dout(1),
            I1 => ram16s_inst_30_dout(1),
            S0 => ad(4)
        );

    mux_inst_135: MUX2
        port map (
            O => mux_o_135,
            I0 => ram16s_inst_32_dout(1),
            I1 => ram16s_inst_34_dout(1),
            S0 => ad(4)
        );

    mux_inst_136: MUX2
        port map (
            O => mux_o_136,
            I0 => ram16s_inst_36_dout(1),
            I1 => ram16s_inst_38_dout(1),
            S0 => ad(4)
        );

    mux_inst_137: MUX2
        port map (
            O => mux_o_137,
            I0 => ram16s_inst_40_dout(1),
            I1 => ram16s_inst_42_dout(1),
            S0 => ad(4)
        );

    mux_inst_138: MUX2
        port map (
            O => mux_o_138,
            I0 => ram16s_inst_44_dout(1),
            I1 => ram16s_inst_46_dout(1),
            S0 => ad(4)
        );

    mux_inst_139: MUX2
        port map (
            O => mux_o_139,
            I0 => ram16s_inst_48_dout(1),
            I1 => ram16s_inst_50_dout(1),
            S0 => ad(4)
        );

    mux_inst_140: MUX2
        port map (
            O => mux_o_140,
            I0 => ram16s_inst_52_dout(1),
            I1 => ram16s_inst_54_dout(1),
            S0 => ad(4)
        );

    mux_inst_141: MUX2
        port map (
            O => mux_o_141,
            I0 => ram16s_inst_56_dout(1),
            I1 => ram16s_inst_58_dout(1),
            S0 => ad(4)
        );

    mux_inst_142: MUX2
        port map (
            O => mux_o_142,
            I0 => ram16s_inst_60_dout(1),
            I1 => ram16s_inst_62_dout(1),
            S0 => ad(4)
        );

    mux_inst_143: MUX2
        port map (
            O => mux_o_143,
            I0 => ram16s_inst_64_dout(1),
            I1 => ram16s_inst_66_dout(1),
            S0 => ad(4)
        );

    mux_inst_144: MUX2
        port map (
            O => mux_o_144,
            I0 => ram16s_inst_68_dout(1),
            I1 => ram16s_inst_70_dout(1),
            S0 => ad(4)
        );

    mux_inst_145: MUX2
        port map (
            O => mux_o_145,
            I0 => ram16s_inst_72_dout(1),
            I1 => ram16s_inst_74_dout(1),
            S0 => ad(4)
        );

    mux_inst_146: MUX2
        port map (
            O => mux_o_146,
            I0 => ram16s_inst_76_dout(1),
            I1 => ram16s_inst_78_dout(1),
            S0 => ad(4)
        );

    mux_inst_147: MUX2
        port map (
            O => mux_o_147,
            I0 => ram16s_inst_80_dout(1),
            I1 => ram16s_inst_82_dout(1),
            S0 => ad(4)
        );

    mux_inst_148: MUX2
        port map (
            O => mux_o_148,
            I0 => ram16s_inst_84_dout(1),
            I1 => ram16s_inst_86_dout(1),
            S0 => ad(4)
        );

    mux_inst_149: MUX2
        port map (
            O => mux_o_149,
            I0 => ram16s_inst_88_dout(1),
            I1 => ram16s_inst_90_dout(1),
            S0 => ad(4)
        );

    mux_inst_150: MUX2
        port map (
            O => mux_o_150,
            I0 => ram16s_inst_92_dout(1),
            I1 => ram16s_inst_94_dout(1),
            S0 => ad(4)
        );

    mux_inst_151: MUX2
        port map (
            O => mux_o_151,
            I0 => ram16s_inst_96_dout(1),
            I1 => ram16s_inst_98_dout(1),
            S0 => ad(4)
        );

    mux_inst_152: MUX2
        port map (
            O => mux_o_152,
            I0 => ram16s_inst_100_dout(1),
            I1 => ram16s_inst_102_dout(1),
            S0 => ad(4)
        );

    mux_inst_153: MUX2
        port map (
            O => mux_o_153,
            I0 => ram16s_inst_104_dout(1),
            I1 => ram16s_inst_106_dout(1),
            S0 => ad(4)
        );

    mux_inst_154: MUX2
        port map (
            O => mux_o_154,
            I0 => ram16s_inst_108_dout(1),
            I1 => ram16s_inst_110_dout(1),
            S0 => ad(4)
        );

    mux_inst_155: MUX2
        port map (
            O => mux_o_155,
            I0 => ram16s_inst_112_dout(1),
            I1 => ram16s_inst_114_dout(1),
            S0 => ad(4)
        );

    mux_inst_156: MUX2
        port map (
            O => mux_o_156,
            I0 => ram16s_inst_116_dout(1),
            I1 => ram16s_inst_118_dout(1),
            S0 => ad(4)
        );

    mux_inst_157: MUX2
        port map (
            O => mux_o_157,
            I0 => ram16s_inst_120_dout(1),
            I1 => ram16s_inst_122_dout(1),
            S0 => ad(4)
        );

    mux_inst_158: MUX2
        port map (
            O => mux_o_158,
            I0 => ram16s_inst_124_dout(1),
            I1 => ram16s_inst_126_dout(1),
            S0 => ad(4)
        );

    mux_inst_159: MUX2
        port map (
            O => mux_o_159,
            I0 => ram16s_inst_128_dout(1),
            I1 => ram16s_inst_130_dout(1),
            S0 => ad(4)
        );

    mux_inst_160: MUX2
        port map (
            O => mux_o_160,
            I0 => ram16s_inst_132_dout(1),
            I1 => ram16s_inst_134_dout(1),
            S0 => ad(4)
        );

    mux_inst_161: MUX2
        port map (
            O => mux_o_161,
            I0 => ram16s_inst_136_dout(1),
            I1 => ram16s_inst_138_dout(1),
            S0 => ad(4)
        );

    mux_inst_162: MUX2
        port map (
            O => mux_o_162,
            I0 => ram16s_inst_140_dout(1),
            I1 => ram16s_inst_142_dout(1),
            S0 => ad(4)
        );

    mux_inst_163: MUX2
        port map (
            O => mux_o_163,
            I0 => ram16s_inst_144_dout(1),
            I1 => ram16s_inst_146_dout(1),
            S0 => ad(4)
        );

    mux_inst_164: MUX2
        port map (
            O => mux_o_164,
            I0 => ram16s_inst_148_dout(1),
            I1 => ram16s_inst_150_dout(1),
            S0 => ad(4)
        );

    mux_inst_165: MUX2
        port map (
            O => mux_o_165,
            I0 => ram16s_inst_152_dout(1),
            I1 => ram16s_inst_154_dout(1),
            S0 => ad(4)
        );

    mux_inst_166: MUX2
        port map (
            O => mux_o_166,
            I0 => ram16s_inst_156_dout(1),
            I1 => ram16s_inst_158_dout(1),
            S0 => ad(4)
        );

    mux_inst_167: MUX2
        port map (
            O => mux_o_167,
            I0 => ram16s_inst_160_dout(1),
            I1 => ram16s_inst_162_dout(1),
            S0 => ad(4)
        );

    mux_inst_168: MUX2
        port map (
            O => mux_o_168,
            I0 => ram16s_inst_164_dout(1),
            I1 => ram16s_inst_166_dout(1),
            S0 => ad(4)
        );

    mux_inst_169: MUX2
        port map (
            O => mux_o_169,
            I0 => ram16s_inst_168_dout(1),
            I1 => ram16s_inst_170_dout(1),
            S0 => ad(4)
        );

    mux_inst_170: MUX2
        port map (
            O => mux_o_170,
            I0 => ram16s_inst_172_dout(1),
            I1 => ram16s_inst_174_dout(1),
            S0 => ad(4)
        );

    mux_inst_171: MUX2
        port map (
            O => mux_o_171,
            I0 => ram16s_inst_176_dout(1),
            I1 => ram16s_inst_178_dout(1),
            S0 => ad(4)
        );

    mux_inst_172: MUX2
        port map (
            O => mux_o_172,
            I0 => ram16s_inst_180_dout(1),
            I1 => ram16s_inst_182_dout(1),
            S0 => ad(4)
        );

    mux_inst_173: MUX2
        port map (
            O => mux_o_173,
            I0 => ram16s_inst_184_dout(1),
            I1 => ram16s_inst_186_dout(1),
            S0 => ad(4)
        );

    mux_inst_174: MUX2
        port map (
            O => mux_o_174,
            I0 => ram16s_inst_188_dout(1),
            I1 => ram16s_inst_190_dout(1),
            S0 => ad(4)
        );

    mux_inst_175: MUX2
        port map (
            O => mux_o_175,
            I0 => ram16s_inst_192_dout(1),
            I1 => ram16s_inst_194_dout(1),
            S0 => ad(4)
        );

    mux_inst_176: MUX2
        port map (
            O => mux_o_176,
            I0 => ram16s_inst_196_dout(1),
            I1 => ram16s_inst_198_dout(1),
            S0 => ad(4)
        );

    mux_inst_177: MUX2
        port map (
            O => mux_o_177,
            I0 => ram16s_inst_200_dout(1),
            I1 => ram16s_inst_202_dout(1),
            S0 => ad(4)
        );

    mux_inst_178: MUX2
        port map (
            O => mux_o_178,
            I0 => ram16s_inst_204_dout(1),
            I1 => ram16s_inst_206_dout(1),
            S0 => ad(4)
        );

    mux_inst_179: MUX2
        port map (
            O => mux_o_179,
            I0 => ram16s_inst_208_dout(1),
            I1 => ram16s_inst_210_dout(1),
            S0 => ad(4)
        );

    mux_inst_180: MUX2
        port map (
            O => mux_o_180,
            I0 => ram16s_inst_212_dout(1),
            I1 => ram16s_inst_214_dout(1),
            S0 => ad(4)
        );

    mux_inst_181: MUX2
        port map (
            O => mux_o_181,
            I0 => ram16s_inst_216_dout(1),
            I1 => ram16s_inst_218_dout(1),
            S0 => ad(4)
        );

    mux_inst_182: MUX2
        port map (
            O => mux_o_182,
            I0 => ram16s_inst_220_dout(1),
            I1 => ram16s_inst_222_dout(1),
            S0 => ad(4)
        );

    mux_inst_183: MUX2
        port map (
            O => mux_o_183,
            I0 => ram16s_inst_224_dout(1),
            I1 => ram16s_inst_226_dout(1),
            S0 => ad(4)
        );

    mux_inst_184: MUX2
        port map (
            O => mux_o_184,
            I0 => ram16s_inst_228_dout(1),
            I1 => ram16s_inst_230_dout(1),
            S0 => ad(4)
        );

    mux_inst_185: MUX2
        port map (
            O => mux_o_185,
            I0 => ram16s_inst_232_dout(1),
            I1 => ram16s_inst_234_dout(1),
            S0 => ad(4)
        );

    mux_inst_186: MUX2
        port map (
            O => mux_o_186,
            I0 => ram16s_inst_236_dout(1),
            I1 => ram16s_inst_238_dout(1),
            S0 => ad(4)
        );

    mux_inst_187: MUX2
        port map (
            O => mux_o_187,
            I0 => ram16s_inst_240_dout(1),
            I1 => ram16s_inst_242_dout(1),
            S0 => ad(4)
        );

    mux_inst_188: MUX2
        port map (
            O => mux_o_188,
            I0 => ram16s_inst_244_dout(1),
            I1 => ram16s_inst_246_dout(1),
            S0 => ad(4)
        );

    mux_inst_189: MUX2
        port map (
            O => mux_o_189,
            I0 => ram16s_inst_248_dout(1),
            I1 => ram16s_inst_250_dout(1),
            S0 => ad(4)
        );

    mux_inst_190: MUX2
        port map (
            O => mux_o_190,
            I0 => ram16s_inst_252_dout(1),
            I1 => ram16s_inst_254_dout(1),
            S0 => ad(4)
        );

    mux_inst_191: MUX2
        port map (
            O => mux_o_191,
            I0 => mux_o_127,
            I1 => mux_o_128,
            S0 => ad(5)
        );

    mux_inst_192: MUX2
        port map (
            O => mux_o_192,
            I0 => mux_o_129,
            I1 => mux_o_130,
            S0 => ad(5)
        );

    mux_inst_193: MUX2
        port map (
            O => mux_o_193,
            I0 => mux_o_131,
            I1 => mux_o_132,
            S0 => ad(5)
        );

    mux_inst_194: MUX2
        port map (
            O => mux_o_194,
            I0 => mux_o_133,
            I1 => mux_o_134,
            S0 => ad(5)
        );

    mux_inst_195: MUX2
        port map (
            O => mux_o_195,
            I0 => mux_o_135,
            I1 => mux_o_136,
            S0 => ad(5)
        );

    mux_inst_196: MUX2
        port map (
            O => mux_o_196,
            I0 => mux_o_137,
            I1 => mux_o_138,
            S0 => ad(5)
        );

    mux_inst_197: MUX2
        port map (
            O => mux_o_197,
            I0 => mux_o_139,
            I1 => mux_o_140,
            S0 => ad(5)
        );

    mux_inst_198: MUX2
        port map (
            O => mux_o_198,
            I0 => mux_o_141,
            I1 => mux_o_142,
            S0 => ad(5)
        );

    mux_inst_199: MUX2
        port map (
            O => mux_o_199,
            I0 => mux_o_143,
            I1 => mux_o_144,
            S0 => ad(5)
        );

    mux_inst_200: MUX2
        port map (
            O => mux_o_200,
            I0 => mux_o_145,
            I1 => mux_o_146,
            S0 => ad(5)
        );

    mux_inst_201: MUX2
        port map (
            O => mux_o_201,
            I0 => mux_o_147,
            I1 => mux_o_148,
            S0 => ad(5)
        );

    mux_inst_202: MUX2
        port map (
            O => mux_o_202,
            I0 => mux_o_149,
            I1 => mux_o_150,
            S0 => ad(5)
        );

    mux_inst_203: MUX2
        port map (
            O => mux_o_203,
            I0 => mux_o_151,
            I1 => mux_o_152,
            S0 => ad(5)
        );

    mux_inst_204: MUX2
        port map (
            O => mux_o_204,
            I0 => mux_o_153,
            I1 => mux_o_154,
            S0 => ad(5)
        );

    mux_inst_205: MUX2
        port map (
            O => mux_o_205,
            I0 => mux_o_155,
            I1 => mux_o_156,
            S0 => ad(5)
        );

    mux_inst_206: MUX2
        port map (
            O => mux_o_206,
            I0 => mux_o_157,
            I1 => mux_o_158,
            S0 => ad(5)
        );

    mux_inst_207: MUX2
        port map (
            O => mux_o_207,
            I0 => mux_o_159,
            I1 => mux_o_160,
            S0 => ad(5)
        );

    mux_inst_208: MUX2
        port map (
            O => mux_o_208,
            I0 => mux_o_161,
            I1 => mux_o_162,
            S0 => ad(5)
        );

    mux_inst_209: MUX2
        port map (
            O => mux_o_209,
            I0 => mux_o_163,
            I1 => mux_o_164,
            S0 => ad(5)
        );

    mux_inst_210: MUX2
        port map (
            O => mux_o_210,
            I0 => mux_o_165,
            I1 => mux_o_166,
            S0 => ad(5)
        );

    mux_inst_211: MUX2
        port map (
            O => mux_o_211,
            I0 => mux_o_167,
            I1 => mux_o_168,
            S0 => ad(5)
        );

    mux_inst_212: MUX2
        port map (
            O => mux_o_212,
            I0 => mux_o_169,
            I1 => mux_o_170,
            S0 => ad(5)
        );

    mux_inst_213: MUX2
        port map (
            O => mux_o_213,
            I0 => mux_o_171,
            I1 => mux_o_172,
            S0 => ad(5)
        );

    mux_inst_214: MUX2
        port map (
            O => mux_o_214,
            I0 => mux_o_173,
            I1 => mux_o_174,
            S0 => ad(5)
        );

    mux_inst_215: MUX2
        port map (
            O => mux_o_215,
            I0 => mux_o_175,
            I1 => mux_o_176,
            S0 => ad(5)
        );

    mux_inst_216: MUX2
        port map (
            O => mux_o_216,
            I0 => mux_o_177,
            I1 => mux_o_178,
            S0 => ad(5)
        );

    mux_inst_217: MUX2
        port map (
            O => mux_o_217,
            I0 => mux_o_179,
            I1 => mux_o_180,
            S0 => ad(5)
        );

    mux_inst_218: MUX2
        port map (
            O => mux_o_218,
            I0 => mux_o_181,
            I1 => mux_o_182,
            S0 => ad(5)
        );

    mux_inst_219: MUX2
        port map (
            O => mux_o_219,
            I0 => mux_o_183,
            I1 => mux_o_184,
            S0 => ad(5)
        );

    mux_inst_220: MUX2
        port map (
            O => mux_o_220,
            I0 => mux_o_185,
            I1 => mux_o_186,
            S0 => ad(5)
        );

    mux_inst_221: MUX2
        port map (
            O => mux_o_221,
            I0 => mux_o_187,
            I1 => mux_o_188,
            S0 => ad(5)
        );

    mux_inst_222: MUX2
        port map (
            O => mux_o_222,
            I0 => mux_o_189,
            I1 => mux_o_190,
            S0 => ad(5)
        );

    mux_inst_223: MUX2
        port map (
            O => mux_o_223,
            I0 => mux_o_191,
            I1 => mux_o_192,
            S0 => ad(6)
        );

    mux_inst_224: MUX2
        port map (
            O => mux_o_224,
            I0 => mux_o_193,
            I1 => mux_o_194,
            S0 => ad(6)
        );

    mux_inst_225: MUX2
        port map (
            O => mux_o_225,
            I0 => mux_o_195,
            I1 => mux_o_196,
            S0 => ad(6)
        );

    mux_inst_226: MUX2
        port map (
            O => mux_o_226,
            I0 => mux_o_197,
            I1 => mux_o_198,
            S0 => ad(6)
        );

    mux_inst_227: MUX2
        port map (
            O => mux_o_227,
            I0 => mux_o_199,
            I1 => mux_o_200,
            S0 => ad(6)
        );

    mux_inst_228: MUX2
        port map (
            O => mux_o_228,
            I0 => mux_o_201,
            I1 => mux_o_202,
            S0 => ad(6)
        );

    mux_inst_229: MUX2
        port map (
            O => mux_o_229,
            I0 => mux_o_203,
            I1 => mux_o_204,
            S0 => ad(6)
        );

    mux_inst_230: MUX2
        port map (
            O => mux_o_230,
            I0 => mux_o_205,
            I1 => mux_o_206,
            S0 => ad(6)
        );

    mux_inst_231: MUX2
        port map (
            O => mux_o_231,
            I0 => mux_o_207,
            I1 => mux_o_208,
            S0 => ad(6)
        );

    mux_inst_232: MUX2
        port map (
            O => mux_o_232,
            I0 => mux_o_209,
            I1 => mux_o_210,
            S0 => ad(6)
        );

    mux_inst_233: MUX2
        port map (
            O => mux_o_233,
            I0 => mux_o_211,
            I1 => mux_o_212,
            S0 => ad(6)
        );

    mux_inst_234: MUX2
        port map (
            O => mux_o_234,
            I0 => mux_o_213,
            I1 => mux_o_214,
            S0 => ad(6)
        );

    mux_inst_235: MUX2
        port map (
            O => mux_o_235,
            I0 => mux_o_215,
            I1 => mux_o_216,
            S0 => ad(6)
        );

    mux_inst_236: MUX2
        port map (
            O => mux_o_236,
            I0 => mux_o_217,
            I1 => mux_o_218,
            S0 => ad(6)
        );

    mux_inst_237: MUX2
        port map (
            O => mux_o_237,
            I0 => mux_o_219,
            I1 => mux_o_220,
            S0 => ad(6)
        );

    mux_inst_238: MUX2
        port map (
            O => mux_o_238,
            I0 => mux_o_221,
            I1 => mux_o_222,
            S0 => ad(6)
        );

    mux_inst_239: MUX2
        port map (
            O => mux_o_239,
            I0 => mux_o_223,
            I1 => mux_o_224,
            S0 => ad(7)
        );

    mux_inst_240: MUX2
        port map (
            O => mux_o_240,
            I0 => mux_o_225,
            I1 => mux_o_226,
            S0 => ad(7)
        );

    mux_inst_241: MUX2
        port map (
            O => mux_o_241,
            I0 => mux_o_227,
            I1 => mux_o_228,
            S0 => ad(7)
        );

    mux_inst_242: MUX2
        port map (
            O => mux_o_242,
            I0 => mux_o_229,
            I1 => mux_o_230,
            S0 => ad(7)
        );

    mux_inst_243: MUX2
        port map (
            O => mux_o_243,
            I0 => mux_o_231,
            I1 => mux_o_232,
            S0 => ad(7)
        );

    mux_inst_244: MUX2
        port map (
            O => mux_o_244,
            I0 => mux_o_233,
            I1 => mux_o_234,
            S0 => ad(7)
        );

    mux_inst_245: MUX2
        port map (
            O => mux_o_245,
            I0 => mux_o_235,
            I1 => mux_o_236,
            S0 => ad(7)
        );

    mux_inst_246: MUX2
        port map (
            O => mux_o_246,
            I0 => mux_o_237,
            I1 => mux_o_238,
            S0 => ad(7)
        );

    mux_inst_247: MUX2
        port map (
            O => mux_o_247,
            I0 => mux_o_239,
            I1 => mux_o_240,
            S0 => ad(8)
        );

    mux_inst_248: MUX2
        port map (
            O => mux_o_248,
            I0 => mux_o_241,
            I1 => mux_o_242,
            S0 => ad(8)
        );

    mux_inst_249: MUX2
        port map (
            O => mux_o_249,
            I0 => mux_o_243,
            I1 => mux_o_244,
            S0 => ad(8)
        );

    mux_inst_250: MUX2
        port map (
            O => mux_o_250,
            I0 => mux_o_245,
            I1 => mux_o_246,
            S0 => ad(8)
        );

    mux_inst_251: MUX2
        port map (
            O => mux_o_251,
            I0 => mux_o_247,
            I1 => mux_o_248,
            S0 => ad(9)
        );

    mux_inst_252: MUX2
        port map (
            O => mux_o_252,
            I0 => mux_o_249,
            I1 => mux_o_250,
            S0 => ad(9)
        );

    mux_inst_253: MUX2
        port map (
            O => dout(1),
            I0 => mux_o_251,
            I1 => mux_o_252,
            S0 => ad(10)
        );

    mux_inst_254: MUX2
        port map (
            O => mux_o_254,
            I0 => ram16s_inst_0_dout(2),
            I1 => ram16s_inst_2_dout(2),
            S0 => ad(4)
        );

    mux_inst_255: MUX2
        port map (
            O => mux_o_255,
            I0 => ram16s_inst_4_dout(2),
            I1 => ram16s_inst_6_dout(2),
            S0 => ad(4)
        );

    mux_inst_256: MUX2
        port map (
            O => mux_o_256,
            I0 => ram16s_inst_8_dout(2),
            I1 => ram16s_inst_10_dout(2),
            S0 => ad(4)
        );

    mux_inst_257: MUX2
        port map (
            O => mux_o_257,
            I0 => ram16s_inst_12_dout(2),
            I1 => ram16s_inst_14_dout(2),
            S0 => ad(4)
        );

    mux_inst_258: MUX2
        port map (
            O => mux_o_258,
            I0 => ram16s_inst_16_dout(2),
            I1 => ram16s_inst_18_dout(2),
            S0 => ad(4)
        );

    mux_inst_259: MUX2
        port map (
            O => mux_o_259,
            I0 => ram16s_inst_20_dout(2),
            I1 => ram16s_inst_22_dout(2),
            S0 => ad(4)
        );

    mux_inst_260: MUX2
        port map (
            O => mux_o_260,
            I0 => ram16s_inst_24_dout(2),
            I1 => ram16s_inst_26_dout(2),
            S0 => ad(4)
        );

    mux_inst_261: MUX2
        port map (
            O => mux_o_261,
            I0 => ram16s_inst_28_dout(2),
            I1 => ram16s_inst_30_dout(2),
            S0 => ad(4)
        );

    mux_inst_262: MUX2
        port map (
            O => mux_o_262,
            I0 => ram16s_inst_32_dout(2),
            I1 => ram16s_inst_34_dout(2),
            S0 => ad(4)
        );

    mux_inst_263: MUX2
        port map (
            O => mux_o_263,
            I0 => ram16s_inst_36_dout(2),
            I1 => ram16s_inst_38_dout(2),
            S0 => ad(4)
        );

    mux_inst_264: MUX2
        port map (
            O => mux_o_264,
            I0 => ram16s_inst_40_dout(2),
            I1 => ram16s_inst_42_dout(2),
            S0 => ad(4)
        );

    mux_inst_265: MUX2
        port map (
            O => mux_o_265,
            I0 => ram16s_inst_44_dout(2),
            I1 => ram16s_inst_46_dout(2),
            S0 => ad(4)
        );

    mux_inst_266: MUX2
        port map (
            O => mux_o_266,
            I0 => ram16s_inst_48_dout(2),
            I1 => ram16s_inst_50_dout(2),
            S0 => ad(4)
        );

    mux_inst_267: MUX2
        port map (
            O => mux_o_267,
            I0 => ram16s_inst_52_dout(2),
            I1 => ram16s_inst_54_dout(2),
            S0 => ad(4)
        );

    mux_inst_268: MUX2
        port map (
            O => mux_o_268,
            I0 => ram16s_inst_56_dout(2),
            I1 => ram16s_inst_58_dout(2),
            S0 => ad(4)
        );

    mux_inst_269: MUX2
        port map (
            O => mux_o_269,
            I0 => ram16s_inst_60_dout(2),
            I1 => ram16s_inst_62_dout(2),
            S0 => ad(4)
        );

    mux_inst_270: MUX2
        port map (
            O => mux_o_270,
            I0 => ram16s_inst_64_dout(2),
            I1 => ram16s_inst_66_dout(2),
            S0 => ad(4)
        );

    mux_inst_271: MUX2
        port map (
            O => mux_o_271,
            I0 => ram16s_inst_68_dout(2),
            I1 => ram16s_inst_70_dout(2),
            S0 => ad(4)
        );

    mux_inst_272: MUX2
        port map (
            O => mux_o_272,
            I0 => ram16s_inst_72_dout(2),
            I1 => ram16s_inst_74_dout(2),
            S0 => ad(4)
        );

    mux_inst_273: MUX2
        port map (
            O => mux_o_273,
            I0 => ram16s_inst_76_dout(2),
            I1 => ram16s_inst_78_dout(2),
            S0 => ad(4)
        );

    mux_inst_274: MUX2
        port map (
            O => mux_o_274,
            I0 => ram16s_inst_80_dout(2),
            I1 => ram16s_inst_82_dout(2),
            S0 => ad(4)
        );

    mux_inst_275: MUX2
        port map (
            O => mux_o_275,
            I0 => ram16s_inst_84_dout(2),
            I1 => ram16s_inst_86_dout(2),
            S0 => ad(4)
        );

    mux_inst_276: MUX2
        port map (
            O => mux_o_276,
            I0 => ram16s_inst_88_dout(2),
            I1 => ram16s_inst_90_dout(2),
            S0 => ad(4)
        );

    mux_inst_277: MUX2
        port map (
            O => mux_o_277,
            I0 => ram16s_inst_92_dout(2),
            I1 => ram16s_inst_94_dout(2),
            S0 => ad(4)
        );

    mux_inst_278: MUX2
        port map (
            O => mux_o_278,
            I0 => ram16s_inst_96_dout(2),
            I1 => ram16s_inst_98_dout(2),
            S0 => ad(4)
        );

    mux_inst_279: MUX2
        port map (
            O => mux_o_279,
            I0 => ram16s_inst_100_dout(2),
            I1 => ram16s_inst_102_dout(2),
            S0 => ad(4)
        );

    mux_inst_280: MUX2
        port map (
            O => mux_o_280,
            I0 => ram16s_inst_104_dout(2),
            I1 => ram16s_inst_106_dout(2),
            S0 => ad(4)
        );

    mux_inst_281: MUX2
        port map (
            O => mux_o_281,
            I0 => ram16s_inst_108_dout(2),
            I1 => ram16s_inst_110_dout(2),
            S0 => ad(4)
        );

    mux_inst_282: MUX2
        port map (
            O => mux_o_282,
            I0 => ram16s_inst_112_dout(2),
            I1 => ram16s_inst_114_dout(2),
            S0 => ad(4)
        );

    mux_inst_283: MUX2
        port map (
            O => mux_o_283,
            I0 => ram16s_inst_116_dout(2),
            I1 => ram16s_inst_118_dout(2),
            S0 => ad(4)
        );

    mux_inst_284: MUX2
        port map (
            O => mux_o_284,
            I0 => ram16s_inst_120_dout(2),
            I1 => ram16s_inst_122_dout(2),
            S0 => ad(4)
        );

    mux_inst_285: MUX2
        port map (
            O => mux_o_285,
            I0 => ram16s_inst_124_dout(2),
            I1 => ram16s_inst_126_dout(2),
            S0 => ad(4)
        );

    mux_inst_286: MUX2
        port map (
            O => mux_o_286,
            I0 => ram16s_inst_128_dout(2),
            I1 => ram16s_inst_130_dout(2),
            S0 => ad(4)
        );

    mux_inst_287: MUX2
        port map (
            O => mux_o_287,
            I0 => ram16s_inst_132_dout(2),
            I1 => ram16s_inst_134_dout(2),
            S0 => ad(4)
        );

    mux_inst_288: MUX2
        port map (
            O => mux_o_288,
            I0 => ram16s_inst_136_dout(2),
            I1 => ram16s_inst_138_dout(2),
            S0 => ad(4)
        );

    mux_inst_289: MUX2
        port map (
            O => mux_o_289,
            I0 => ram16s_inst_140_dout(2),
            I1 => ram16s_inst_142_dout(2),
            S0 => ad(4)
        );

    mux_inst_290: MUX2
        port map (
            O => mux_o_290,
            I0 => ram16s_inst_144_dout(2),
            I1 => ram16s_inst_146_dout(2),
            S0 => ad(4)
        );

    mux_inst_291: MUX2
        port map (
            O => mux_o_291,
            I0 => ram16s_inst_148_dout(2),
            I1 => ram16s_inst_150_dout(2),
            S0 => ad(4)
        );

    mux_inst_292: MUX2
        port map (
            O => mux_o_292,
            I0 => ram16s_inst_152_dout(2),
            I1 => ram16s_inst_154_dout(2),
            S0 => ad(4)
        );

    mux_inst_293: MUX2
        port map (
            O => mux_o_293,
            I0 => ram16s_inst_156_dout(2),
            I1 => ram16s_inst_158_dout(2),
            S0 => ad(4)
        );

    mux_inst_294: MUX2
        port map (
            O => mux_o_294,
            I0 => ram16s_inst_160_dout(2),
            I1 => ram16s_inst_162_dout(2),
            S0 => ad(4)
        );

    mux_inst_295: MUX2
        port map (
            O => mux_o_295,
            I0 => ram16s_inst_164_dout(2),
            I1 => ram16s_inst_166_dout(2),
            S0 => ad(4)
        );

    mux_inst_296: MUX2
        port map (
            O => mux_o_296,
            I0 => ram16s_inst_168_dout(2),
            I1 => ram16s_inst_170_dout(2),
            S0 => ad(4)
        );

    mux_inst_297: MUX2
        port map (
            O => mux_o_297,
            I0 => ram16s_inst_172_dout(2),
            I1 => ram16s_inst_174_dout(2),
            S0 => ad(4)
        );

    mux_inst_298: MUX2
        port map (
            O => mux_o_298,
            I0 => ram16s_inst_176_dout(2),
            I1 => ram16s_inst_178_dout(2),
            S0 => ad(4)
        );

    mux_inst_299: MUX2
        port map (
            O => mux_o_299,
            I0 => ram16s_inst_180_dout(2),
            I1 => ram16s_inst_182_dout(2),
            S0 => ad(4)
        );

    mux_inst_300: MUX2
        port map (
            O => mux_o_300,
            I0 => ram16s_inst_184_dout(2),
            I1 => ram16s_inst_186_dout(2),
            S0 => ad(4)
        );

    mux_inst_301: MUX2
        port map (
            O => mux_o_301,
            I0 => ram16s_inst_188_dout(2),
            I1 => ram16s_inst_190_dout(2),
            S0 => ad(4)
        );

    mux_inst_302: MUX2
        port map (
            O => mux_o_302,
            I0 => ram16s_inst_192_dout(2),
            I1 => ram16s_inst_194_dout(2),
            S0 => ad(4)
        );

    mux_inst_303: MUX2
        port map (
            O => mux_o_303,
            I0 => ram16s_inst_196_dout(2),
            I1 => ram16s_inst_198_dout(2),
            S0 => ad(4)
        );

    mux_inst_304: MUX2
        port map (
            O => mux_o_304,
            I0 => ram16s_inst_200_dout(2),
            I1 => ram16s_inst_202_dout(2),
            S0 => ad(4)
        );

    mux_inst_305: MUX2
        port map (
            O => mux_o_305,
            I0 => ram16s_inst_204_dout(2),
            I1 => ram16s_inst_206_dout(2),
            S0 => ad(4)
        );

    mux_inst_306: MUX2
        port map (
            O => mux_o_306,
            I0 => ram16s_inst_208_dout(2),
            I1 => ram16s_inst_210_dout(2),
            S0 => ad(4)
        );

    mux_inst_307: MUX2
        port map (
            O => mux_o_307,
            I0 => ram16s_inst_212_dout(2),
            I1 => ram16s_inst_214_dout(2),
            S0 => ad(4)
        );

    mux_inst_308: MUX2
        port map (
            O => mux_o_308,
            I0 => ram16s_inst_216_dout(2),
            I1 => ram16s_inst_218_dout(2),
            S0 => ad(4)
        );

    mux_inst_309: MUX2
        port map (
            O => mux_o_309,
            I0 => ram16s_inst_220_dout(2),
            I1 => ram16s_inst_222_dout(2),
            S0 => ad(4)
        );

    mux_inst_310: MUX2
        port map (
            O => mux_o_310,
            I0 => ram16s_inst_224_dout(2),
            I1 => ram16s_inst_226_dout(2),
            S0 => ad(4)
        );

    mux_inst_311: MUX2
        port map (
            O => mux_o_311,
            I0 => ram16s_inst_228_dout(2),
            I1 => ram16s_inst_230_dout(2),
            S0 => ad(4)
        );

    mux_inst_312: MUX2
        port map (
            O => mux_o_312,
            I0 => ram16s_inst_232_dout(2),
            I1 => ram16s_inst_234_dout(2),
            S0 => ad(4)
        );

    mux_inst_313: MUX2
        port map (
            O => mux_o_313,
            I0 => ram16s_inst_236_dout(2),
            I1 => ram16s_inst_238_dout(2),
            S0 => ad(4)
        );

    mux_inst_314: MUX2
        port map (
            O => mux_o_314,
            I0 => ram16s_inst_240_dout(2),
            I1 => ram16s_inst_242_dout(2),
            S0 => ad(4)
        );

    mux_inst_315: MUX2
        port map (
            O => mux_o_315,
            I0 => ram16s_inst_244_dout(2),
            I1 => ram16s_inst_246_dout(2),
            S0 => ad(4)
        );

    mux_inst_316: MUX2
        port map (
            O => mux_o_316,
            I0 => ram16s_inst_248_dout(2),
            I1 => ram16s_inst_250_dout(2),
            S0 => ad(4)
        );

    mux_inst_317: MUX2
        port map (
            O => mux_o_317,
            I0 => ram16s_inst_252_dout(2),
            I1 => ram16s_inst_254_dout(2),
            S0 => ad(4)
        );

    mux_inst_318: MUX2
        port map (
            O => mux_o_318,
            I0 => mux_o_254,
            I1 => mux_o_255,
            S0 => ad(5)
        );

    mux_inst_319: MUX2
        port map (
            O => mux_o_319,
            I0 => mux_o_256,
            I1 => mux_o_257,
            S0 => ad(5)
        );

    mux_inst_320: MUX2
        port map (
            O => mux_o_320,
            I0 => mux_o_258,
            I1 => mux_o_259,
            S0 => ad(5)
        );

    mux_inst_321: MUX2
        port map (
            O => mux_o_321,
            I0 => mux_o_260,
            I1 => mux_o_261,
            S0 => ad(5)
        );

    mux_inst_322: MUX2
        port map (
            O => mux_o_322,
            I0 => mux_o_262,
            I1 => mux_o_263,
            S0 => ad(5)
        );

    mux_inst_323: MUX2
        port map (
            O => mux_o_323,
            I0 => mux_o_264,
            I1 => mux_o_265,
            S0 => ad(5)
        );

    mux_inst_324: MUX2
        port map (
            O => mux_o_324,
            I0 => mux_o_266,
            I1 => mux_o_267,
            S0 => ad(5)
        );

    mux_inst_325: MUX2
        port map (
            O => mux_o_325,
            I0 => mux_o_268,
            I1 => mux_o_269,
            S0 => ad(5)
        );

    mux_inst_326: MUX2
        port map (
            O => mux_o_326,
            I0 => mux_o_270,
            I1 => mux_o_271,
            S0 => ad(5)
        );

    mux_inst_327: MUX2
        port map (
            O => mux_o_327,
            I0 => mux_o_272,
            I1 => mux_o_273,
            S0 => ad(5)
        );

    mux_inst_328: MUX2
        port map (
            O => mux_o_328,
            I0 => mux_o_274,
            I1 => mux_o_275,
            S0 => ad(5)
        );

    mux_inst_329: MUX2
        port map (
            O => mux_o_329,
            I0 => mux_o_276,
            I1 => mux_o_277,
            S0 => ad(5)
        );

    mux_inst_330: MUX2
        port map (
            O => mux_o_330,
            I0 => mux_o_278,
            I1 => mux_o_279,
            S0 => ad(5)
        );

    mux_inst_331: MUX2
        port map (
            O => mux_o_331,
            I0 => mux_o_280,
            I1 => mux_o_281,
            S0 => ad(5)
        );

    mux_inst_332: MUX2
        port map (
            O => mux_o_332,
            I0 => mux_o_282,
            I1 => mux_o_283,
            S0 => ad(5)
        );

    mux_inst_333: MUX2
        port map (
            O => mux_o_333,
            I0 => mux_o_284,
            I1 => mux_o_285,
            S0 => ad(5)
        );

    mux_inst_334: MUX2
        port map (
            O => mux_o_334,
            I0 => mux_o_286,
            I1 => mux_o_287,
            S0 => ad(5)
        );

    mux_inst_335: MUX2
        port map (
            O => mux_o_335,
            I0 => mux_o_288,
            I1 => mux_o_289,
            S0 => ad(5)
        );

    mux_inst_336: MUX2
        port map (
            O => mux_o_336,
            I0 => mux_o_290,
            I1 => mux_o_291,
            S0 => ad(5)
        );

    mux_inst_337: MUX2
        port map (
            O => mux_o_337,
            I0 => mux_o_292,
            I1 => mux_o_293,
            S0 => ad(5)
        );

    mux_inst_338: MUX2
        port map (
            O => mux_o_338,
            I0 => mux_o_294,
            I1 => mux_o_295,
            S0 => ad(5)
        );

    mux_inst_339: MUX2
        port map (
            O => mux_o_339,
            I0 => mux_o_296,
            I1 => mux_o_297,
            S0 => ad(5)
        );

    mux_inst_340: MUX2
        port map (
            O => mux_o_340,
            I0 => mux_o_298,
            I1 => mux_o_299,
            S0 => ad(5)
        );

    mux_inst_341: MUX2
        port map (
            O => mux_o_341,
            I0 => mux_o_300,
            I1 => mux_o_301,
            S0 => ad(5)
        );

    mux_inst_342: MUX2
        port map (
            O => mux_o_342,
            I0 => mux_o_302,
            I1 => mux_o_303,
            S0 => ad(5)
        );

    mux_inst_343: MUX2
        port map (
            O => mux_o_343,
            I0 => mux_o_304,
            I1 => mux_o_305,
            S0 => ad(5)
        );

    mux_inst_344: MUX2
        port map (
            O => mux_o_344,
            I0 => mux_o_306,
            I1 => mux_o_307,
            S0 => ad(5)
        );

    mux_inst_345: MUX2
        port map (
            O => mux_o_345,
            I0 => mux_o_308,
            I1 => mux_o_309,
            S0 => ad(5)
        );

    mux_inst_346: MUX2
        port map (
            O => mux_o_346,
            I0 => mux_o_310,
            I1 => mux_o_311,
            S0 => ad(5)
        );

    mux_inst_347: MUX2
        port map (
            O => mux_o_347,
            I0 => mux_o_312,
            I1 => mux_o_313,
            S0 => ad(5)
        );

    mux_inst_348: MUX2
        port map (
            O => mux_o_348,
            I0 => mux_o_314,
            I1 => mux_o_315,
            S0 => ad(5)
        );

    mux_inst_349: MUX2
        port map (
            O => mux_o_349,
            I0 => mux_o_316,
            I1 => mux_o_317,
            S0 => ad(5)
        );

    mux_inst_350: MUX2
        port map (
            O => mux_o_350,
            I0 => mux_o_318,
            I1 => mux_o_319,
            S0 => ad(6)
        );

    mux_inst_351: MUX2
        port map (
            O => mux_o_351,
            I0 => mux_o_320,
            I1 => mux_o_321,
            S0 => ad(6)
        );

    mux_inst_352: MUX2
        port map (
            O => mux_o_352,
            I0 => mux_o_322,
            I1 => mux_o_323,
            S0 => ad(6)
        );

    mux_inst_353: MUX2
        port map (
            O => mux_o_353,
            I0 => mux_o_324,
            I1 => mux_o_325,
            S0 => ad(6)
        );

    mux_inst_354: MUX2
        port map (
            O => mux_o_354,
            I0 => mux_o_326,
            I1 => mux_o_327,
            S0 => ad(6)
        );

    mux_inst_355: MUX2
        port map (
            O => mux_o_355,
            I0 => mux_o_328,
            I1 => mux_o_329,
            S0 => ad(6)
        );

    mux_inst_356: MUX2
        port map (
            O => mux_o_356,
            I0 => mux_o_330,
            I1 => mux_o_331,
            S0 => ad(6)
        );

    mux_inst_357: MUX2
        port map (
            O => mux_o_357,
            I0 => mux_o_332,
            I1 => mux_o_333,
            S0 => ad(6)
        );

    mux_inst_358: MUX2
        port map (
            O => mux_o_358,
            I0 => mux_o_334,
            I1 => mux_o_335,
            S0 => ad(6)
        );

    mux_inst_359: MUX2
        port map (
            O => mux_o_359,
            I0 => mux_o_336,
            I1 => mux_o_337,
            S0 => ad(6)
        );

    mux_inst_360: MUX2
        port map (
            O => mux_o_360,
            I0 => mux_o_338,
            I1 => mux_o_339,
            S0 => ad(6)
        );

    mux_inst_361: MUX2
        port map (
            O => mux_o_361,
            I0 => mux_o_340,
            I1 => mux_o_341,
            S0 => ad(6)
        );

    mux_inst_362: MUX2
        port map (
            O => mux_o_362,
            I0 => mux_o_342,
            I1 => mux_o_343,
            S0 => ad(6)
        );

    mux_inst_363: MUX2
        port map (
            O => mux_o_363,
            I0 => mux_o_344,
            I1 => mux_o_345,
            S0 => ad(6)
        );

    mux_inst_364: MUX2
        port map (
            O => mux_o_364,
            I0 => mux_o_346,
            I1 => mux_o_347,
            S0 => ad(6)
        );

    mux_inst_365: MUX2
        port map (
            O => mux_o_365,
            I0 => mux_o_348,
            I1 => mux_o_349,
            S0 => ad(6)
        );

    mux_inst_366: MUX2
        port map (
            O => mux_o_366,
            I0 => mux_o_350,
            I1 => mux_o_351,
            S0 => ad(7)
        );

    mux_inst_367: MUX2
        port map (
            O => mux_o_367,
            I0 => mux_o_352,
            I1 => mux_o_353,
            S0 => ad(7)
        );

    mux_inst_368: MUX2
        port map (
            O => mux_o_368,
            I0 => mux_o_354,
            I1 => mux_o_355,
            S0 => ad(7)
        );

    mux_inst_369: MUX2
        port map (
            O => mux_o_369,
            I0 => mux_o_356,
            I1 => mux_o_357,
            S0 => ad(7)
        );

    mux_inst_370: MUX2
        port map (
            O => mux_o_370,
            I0 => mux_o_358,
            I1 => mux_o_359,
            S0 => ad(7)
        );

    mux_inst_371: MUX2
        port map (
            O => mux_o_371,
            I0 => mux_o_360,
            I1 => mux_o_361,
            S0 => ad(7)
        );

    mux_inst_372: MUX2
        port map (
            O => mux_o_372,
            I0 => mux_o_362,
            I1 => mux_o_363,
            S0 => ad(7)
        );

    mux_inst_373: MUX2
        port map (
            O => mux_o_373,
            I0 => mux_o_364,
            I1 => mux_o_365,
            S0 => ad(7)
        );

    mux_inst_374: MUX2
        port map (
            O => mux_o_374,
            I0 => mux_o_366,
            I1 => mux_o_367,
            S0 => ad(8)
        );

    mux_inst_375: MUX2
        port map (
            O => mux_o_375,
            I0 => mux_o_368,
            I1 => mux_o_369,
            S0 => ad(8)
        );

    mux_inst_376: MUX2
        port map (
            O => mux_o_376,
            I0 => mux_o_370,
            I1 => mux_o_371,
            S0 => ad(8)
        );

    mux_inst_377: MUX2
        port map (
            O => mux_o_377,
            I0 => mux_o_372,
            I1 => mux_o_373,
            S0 => ad(8)
        );

    mux_inst_378: MUX2
        port map (
            O => mux_o_378,
            I0 => mux_o_374,
            I1 => mux_o_375,
            S0 => ad(9)
        );

    mux_inst_379: MUX2
        port map (
            O => mux_o_379,
            I0 => mux_o_376,
            I1 => mux_o_377,
            S0 => ad(9)
        );

    mux_inst_380: MUX2
        port map (
            O => dout(2),
            I0 => mux_o_378,
            I1 => mux_o_379,
            S0 => ad(10)
        );

    mux_inst_381: MUX2
        port map (
            O => mux_o_381,
            I0 => ram16s_inst_0_dout(3),
            I1 => ram16s_inst_2_dout(3),
            S0 => ad(4)
        );

    mux_inst_382: MUX2
        port map (
            O => mux_o_382,
            I0 => ram16s_inst_4_dout(3),
            I1 => ram16s_inst_6_dout(3),
            S0 => ad(4)
        );

    mux_inst_383: MUX2
        port map (
            O => mux_o_383,
            I0 => ram16s_inst_8_dout(3),
            I1 => ram16s_inst_10_dout(3),
            S0 => ad(4)
        );

    mux_inst_384: MUX2
        port map (
            O => mux_o_384,
            I0 => ram16s_inst_12_dout(3),
            I1 => ram16s_inst_14_dout(3),
            S0 => ad(4)
        );

    mux_inst_385: MUX2
        port map (
            O => mux_o_385,
            I0 => ram16s_inst_16_dout(3),
            I1 => ram16s_inst_18_dout(3),
            S0 => ad(4)
        );

    mux_inst_386: MUX2
        port map (
            O => mux_o_386,
            I0 => ram16s_inst_20_dout(3),
            I1 => ram16s_inst_22_dout(3),
            S0 => ad(4)
        );

    mux_inst_387: MUX2
        port map (
            O => mux_o_387,
            I0 => ram16s_inst_24_dout(3),
            I1 => ram16s_inst_26_dout(3),
            S0 => ad(4)
        );

    mux_inst_388: MUX2
        port map (
            O => mux_o_388,
            I0 => ram16s_inst_28_dout(3),
            I1 => ram16s_inst_30_dout(3),
            S0 => ad(4)
        );

    mux_inst_389: MUX2
        port map (
            O => mux_o_389,
            I0 => ram16s_inst_32_dout(3),
            I1 => ram16s_inst_34_dout(3),
            S0 => ad(4)
        );

    mux_inst_390: MUX2
        port map (
            O => mux_o_390,
            I0 => ram16s_inst_36_dout(3),
            I1 => ram16s_inst_38_dout(3),
            S0 => ad(4)
        );

    mux_inst_391: MUX2
        port map (
            O => mux_o_391,
            I0 => ram16s_inst_40_dout(3),
            I1 => ram16s_inst_42_dout(3),
            S0 => ad(4)
        );

    mux_inst_392: MUX2
        port map (
            O => mux_o_392,
            I0 => ram16s_inst_44_dout(3),
            I1 => ram16s_inst_46_dout(3),
            S0 => ad(4)
        );

    mux_inst_393: MUX2
        port map (
            O => mux_o_393,
            I0 => ram16s_inst_48_dout(3),
            I1 => ram16s_inst_50_dout(3),
            S0 => ad(4)
        );

    mux_inst_394: MUX2
        port map (
            O => mux_o_394,
            I0 => ram16s_inst_52_dout(3),
            I1 => ram16s_inst_54_dout(3),
            S0 => ad(4)
        );

    mux_inst_395: MUX2
        port map (
            O => mux_o_395,
            I0 => ram16s_inst_56_dout(3),
            I1 => ram16s_inst_58_dout(3),
            S0 => ad(4)
        );

    mux_inst_396: MUX2
        port map (
            O => mux_o_396,
            I0 => ram16s_inst_60_dout(3),
            I1 => ram16s_inst_62_dout(3),
            S0 => ad(4)
        );

    mux_inst_397: MUX2
        port map (
            O => mux_o_397,
            I0 => ram16s_inst_64_dout(3),
            I1 => ram16s_inst_66_dout(3),
            S0 => ad(4)
        );

    mux_inst_398: MUX2
        port map (
            O => mux_o_398,
            I0 => ram16s_inst_68_dout(3),
            I1 => ram16s_inst_70_dout(3),
            S0 => ad(4)
        );

    mux_inst_399: MUX2
        port map (
            O => mux_o_399,
            I0 => ram16s_inst_72_dout(3),
            I1 => ram16s_inst_74_dout(3),
            S0 => ad(4)
        );

    mux_inst_400: MUX2
        port map (
            O => mux_o_400,
            I0 => ram16s_inst_76_dout(3),
            I1 => ram16s_inst_78_dout(3),
            S0 => ad(4)
        );

    mux_inst_401: MUX2
        port map (
            O => mux_o_401,
            I0 => ram16s_inst_80_dout(3),
            I1 => ram16s_inst_82_dout(3),
            S0 => ad(4)
        );

    mux_inst_402: MUX2
        port map (
            O => mux_o_402,
            I0 => ram16s_inst_84_dout(3),
            I1 => ram16s_inst_86_dout(3),
            S0 => ad(4)
        );

    mux_inst_403: MUX2
        port map (
            O => mux_o_403,
            I0 => ram16s_inst_88_dout(3),
            I1 => ram16s_inst_90_dout(3),
            S0 => ad(4)
        );

    mux_inst_404: MUX2
        port map (
            O => mux_o_404,
            I0 => ram16s_inst_92_dout(3),
            I1 => ram16s_inst_94_dout(3),
            S0 => ad(4)
        );

    mux_inst_405: MUX2
        port map (
            O => mux_o_405,
            I0 => ram16s_inst_96_dout(3),
            I1 => ram16s_inst_98_dout(3),
            S0 => ad(4)
        );

    mux_inst_406: MUX2
        port map (
            O => mux_o_406,
            I0 => ram16s_inst_100_dout(3),
            I1 => ram16s_inst_102_dout(3),
            S0 => ad(4)
        );

    mux_inst_407: MUX2
        port map (
            O => mux_o_407,
            I0 => ram16s_inst_104_dout(3),
            I1 => ram16s_inst_106_dout(3),
            S0 => ad(4)
        );

    mux_inst_408: MUX2
        port map (
            O => mux_o_408,
            I0 => ram16s_inst_108_dout(3),
            I1 => ram16s_inst_110_dout(3),
            S0 => ad(4)
        );

    mux_inst_409: MUX2
        port map (
            O => mux_o_409,
            I0 => ram16s_inst_112_dout(3),
            I1 => ram16s_inst_114_dout(3),
            S0 => ad(4)
        );

    mux_inst_410: MUX2
        port map (
            O => mux_o_410,
            I0 => ram16s_inst_116_dout(3),
            I1 => ram16s_inst_118_dout(3),
            S0 => ad(4)
        );

    mux_inst_411: MUX2
        port map (
            O => mux_o_411,
            I0 => ram16s_inst_120_dout(3),
            I1 => ram16s_inst_122_dout(3),
            S0 => ad(4)
        );

    mux_inst_412: MUX2
        port map (
            O => mux_o_412,
            I0 => ram16s_inst_124_dout(3),
            I1 => ram16s_inst_126_dout(3),
            S0 => ad(4)
        );

    mux_inst_413: MUX2
        port map (
            O => mux_o_413,
            I0 => ram16s_inst_128_dout(3),
            I1 => ram16s_inst_130_dout(3),
            S0 => ad(4)
        );

    mux_inst_414: MUX2
        port map (
            O => mux_o_414,
            I0 => ram16s_inst_132_dout(3),
            I1 => ram16s_inst_134_dout(3),
            S0 => ad(4)
        );

    mux_inst_415: MUX2
        port map (
            O => mux_o_415,
            I0 => ram16s_inst_136_dout(3),
            I1 => ram16s_inst_138_dout(3),
            S0 => ad(4)
        );

    mux_inst_416: MUX2
        port map (
            O => mux_o_416,
            I0 => ram16s_inst_140_dout(3),
            I1 => ram16s_inst_142_dout(3),
            S0 => ad(4)
        );

    mux_inst_417: MUX2
        port map (
            O => mux_o_417,
            I0 => ram16s_inst_144_dout(3),
            I1 => ram16s_inst_146_dout(3),
            S0 => ad(4)
        );

    mux_inst_418: MUX2
        port map (
            O => mux_o_418,
            I0 => ram16s_inst_148_dout(3),
            I1 => ram16s_inst_150_dout(3),
            S0 => ad(4)
        );

    mux_inst_419: MUX2
        port map (
            O => mux_o_419,
            I0 => ram16s_inst_152_dout(3),
            I1 => ram16s_inst_154_dout(3),
            S0 => ad(4)
        );

    mux_inst_420: MUX2
        port map (
            O => mux_o_420,
            I0 => ram16s_inst_156_dout(3),
            I1 => ram16s_inst_158_dout(3),
            S0 => ad(4)
        );

    mux_inst_421: MUX2
        port map (
            O => mux_o_421,
            I0 => ram16s_inst_160_dout(3),
            I1 => ram16s_inst_162_dout(3),
            S0 => ad(4)
        );

    mux_inst_422: MUX2
        port map (
            O => mux_o_422,
            I0 => ram16s_inst_164_dout(3),
            I1 => ram16s_inst_166_dout(3),
            S0 => ad(4)
        );

    mux_inst_423: MUX2
        port map (
            O => mux_o_423,
            I0 => ram16s_inst_168_dout(3),
            I1 => ram16s_inst_170_dout(3),
            S0 => ad(4)
        );

    mux_inst_424: MUX2
        port map (
            O => mux_o_424,
            I0 => ram16s_inst_172_dout(3),
            I1 => ram16s_inst_174_dout(3),
            S0 => ad(4)
        );

    mux_inst_425: MUX2
        port map (
            O => mux_o_425,
            I0 => ram16s_inst_176_dout(3),
            I1 => ram16s_inst_178_dout(3),
            S0 => ad(4)
        );

    mux_inst_426: MUX2
        port map (
            O => mux_o_426,
            I0 => ram16s_inst_180_dout(3),
            I1 => ram16s_inst_182_dout(3),
            S0 => ad(4)
        );

    mux_inst_427: MUX2
        port map (
            O => mux_o_427,
            I0 => ram16s_inst_184_dout(3),
            I1 => ram16s_inst_186_dout(3),
            S0 => ad(4)
        );

    mux_inst_428: MUX2
        port map (
            O => mux_o_428,
            I0 => ram16s_inst_188_dout(3),
            I1 => ram16s_inst_190_dout(3),
            S0 => ad(4)
        );

    mux_inst_429: MUX2
        port map (
            O => mux_o_429,
            I0 => ram16s_inst_192_dout(3),
            I1 => ram16s_inst_194_dout(3),
            S0 => ad(4)
        );

    mux_inst_430: MUX2
        port map (
            O => mux_o_430,
            I0 => ram16s_inst_196_dout(3),
            I1 => ram16s_inst_198_dout(3),
            S0 => ad(4)
        );

    mux_inst_431: MUX2
        port map (
            O => mux_o_431,
            I0 => ram16s_inst_200_dout(3),
            I1 => ram16s_inst_202_dout(3),
            S0 => ad(4)
        );

    mux_inst_432: MUX2
        port map (
            O => mux_o_432,
            I0 => ram16s_inst_204_dout(3),
            I1 => ram16s_inst_206_dout(3),
            S0 => ad(4)
        );

    mux_inst_433: MUX2
        port map (
            O => mux_o_433,
            I0 => ram16s_inst_208_dout(3),
            I1 => ram16s_inst_210_dout(3),
            S0 => ad(4)
        );

    mux_inst_434: MUX2
        port map (
            O => mux_o_434,
            I0 => ram16s_inst_212_dout(3),
            I1 => ram16s_inst_214_dout(3),
            S0 => ad(4)
        );

    mux_inst_435: MUX2
        port map (
            O => mux_o_435,
            I0 => ram16s_inst_216_dout(3),
            I1 => ram16s_inst_218_dout(3),
            S0 => ad(4)
        );

    mux_inst_436: MUX2
        port map (
            O => mux_o_436,
            I0 => ram16s_inst_220_dout(3),
            I1 => ram16s_inst_222_dout(3),
            S0 => ad(4)
        );

    mux_inst_437: MUX2
        port map (
            O => mux_o_437,
            I0 => ram16s_inst_224_dout(3),
            I1 => ram16s_inst_226_dout(3),
            S0 => ad(4)
        );

    mux_inst_438: MUX2
        port map (
            O => mux_o_438,
            I0 => ram16s_inst_228_dout(3),
            I1 => ram16s_inst_230_dout(3),
            S0 => ad(4)
        );

    mux_inst_439: MUX2
        port map (
            O => mux_o_439,
            I0 => ram16s_inst_232_dout(3),
            I1 => ram16s_inst_234_dout(3),
            S0 => ad(4)
        );

    mux_inst_440: MUX2
        port map (
            O => mux_o_440,
            I0 => ram16s_inst_236_dout(3),
            I1 => ram16s_inst_238_dout(3),
            S0 => ad(4)
        );

    mux_inst_441: MUX2
        port map (
            O => mux_o_441,
            I0 => ram16s_inst_240_dout(3),
            I1 => ram16s_inst_242_dout(3),
            S0 => ad(4)
        );

    mux_inst_442: MUX2
        port map (
            O => mux_o_442,
            I0 => ram16s_inst_244_dout(3),
            I1 => ram16s_inst_246_dout(3),
            S0 => ad(4)
        );

    mux_inst_443: MUX2
        port map (
            O => mux_o_443,
            I0 => ram16s_inst_248_dout(3),
            I1 => ram16s_inst_250_dout(3),
            S0 => ad(4)
        );

    mux_inst_444: MUX2
        port map (
            O => mux_o_444,
            I0 => ram16s_inst_252_dout(3),
            I1 => ram16s_inst_254_dout(3),
            S0 => ad(4)
        );

    mux_inst_445: MUX2
        port map (
            O => mux_o_445,
            I0 => mux_o_381,
            I1 => mux_o_382,
            S0 => ad(5)
        );

    mux_inst_446: MUX2
        port map (
            O => mux_o_446,
            I0 => mux_o_383,
            I1 => mux_o_384,
            S0 => ad(5)
        );

    mux_inst_447: MUX2
        port map (
            O => mux_o_447,
            I0 => mux_o_385,
            I1 => mux_o_386,
            S0 => ad(5)
        );

    mux_inst_448: MUX2
        port map (
            O => mux_o_448,
            I0 => mux_o_387,
            I1 => mux_o_388,
            S0 => ad(5)
        );

    mux_inst_449: MUX2
        port map (
            O => mux_o_449,
            I0 => mux_o_389,
            I1 => mux_o_390,
            S0 => ad(5)
        );

    mux_inst_450: MUX2
        port map (
            O => mux_o_450,
            I0 => mux_o_391,
            I1 => mux_o_392,
            S0 => ad(5)
        );

    mux_inst_451: MUX2
        port map (
            O => mux_o_451,
            I0 => mux_o_393,
            I1 => mux_o_394,
            S0 => ad(5)
        );

    mux_inst_452: MUX2
        port map (
            O => mux_o_452,
            I0 => mux_o_395,
            I1 => mux_o_396,
            S0 => ad(5)
        );

    mux_inst_453: MUX2
        port map (
            O => mux_o_453,
            I0 => mux_o_397,
            I1 => mux_o_398,
            S0 => ad(5)
        );

    mux_inst_454: MUX2
        port map (
            O => mux_o_454,
            I0 => mux_o_399,
            I1 => mux_o_400,
            S0 => ad(5)
        );

    mux_inst_455: MUX2
        port map (
            O => mux_o_455,
            I0 => mux_o_401,
            I1 => mux_o_402,
            S0 => ad(5)
        );

    mux_inst_456: MUX2
        port map (
            O => mux_o_456,
            I0 => mux_o_403,
            I1 => mux_o_404,
            S0 => ad(5)
        );

    mux_inst_457: MUX2
        port map (
            O => mux_o_457,
            I0 => mux_o_405,
            I1 => mux_o_406,
            S0 => ad(5)
        );

    mux_inst_458: MUX2
        port map (
            O => mux_o_458,
            I0 => mux_o_407,
            I1 => mux_o_408,
            S0 => ad(5)
        );

    mux_inst_459: MUX2
        port map (
            O => mux_o_459,
            I0 => mux_o_409,
            I1 => mux_o_410,
            S0 => ad(5)
        );

    mux_inst_460: MUX2
        port map (
            O => mux_o_460,
            I0 => mux_o_411,
            I1 => mux_o_412,
            S0 => ad(5)
        );

    mux_inst_461: MUX2
        port map (
            O => mux_o_461,
            I0 => mux_o_413,
            I1 => mux_o_414,
            S0 => ad(5)
        );

    mux_inst_462: MUX2
        port map (
            O => mux_o_462,
            I0 => mux_o_415,
            I1 => mux_o_416,
            S0 => ad(5)
        );

    mux_inst_463: MUX2
        port map (
            O => mux_o_463,
            I0 => mux_o_417,
            I1 => mux_o_418,
            S0 => ad(5)
        );

    mux_inst_464: MUX2
        port map (
            O => mux_o_464,
            I0 => mux_o_419,
            I1 => mux_o_420,
            S0 => ad(5)
        );

    mux_inst_465: MUX2
        port map (
            O => mux_o_465,
            I0 => mux_o_421,
            I1 => mux_o_422,
            S0 => ad(5)
        );

    mux_inst_466: MUX2
        port map (
            O => mux_o_466,
            I0 => mux_o_423,
            I1 => mux_o_424,
            S0 => ad(5)
        );

    mux_inst_467: MUX2
        port map (
            O => mux_o_467,
            I0 => mux_o_425,
            I1 => mux_o_426,
            S0 => ad(5)
        );

    mux_inst_468: MUX2
        port map (
            O => mux_o_468,
            I0 => mux_o_427,
            I1 => mux_o_428,
            S0 => ad(5)
        );

    mux_inst_469: MUX2
        port map (
            O => mux_o_469,
            I0 => mux_o_429,
            I1 => mux_o_430,
            S0 => ad(5)
        );

    mux_inst_470: MUX2
        port map (
            O => mux_o_470,
            I0 => mux_o_431,
            I1 => mux_o_432,
            S0 => ad(5)
        );

    mux_inst_471: MUX2
        port map (
            O => mux_o_471,
            I0 => mux_o_433,
            I1 => mux_o_434,
            S0 => ad(5)
        );

    mux_inst_472: MUX2
        port map (
            O => mux_o_472,
            I0 => mux_o_435,
            I1 => mux_o_436,
            S0 => ad(5)
        );

    mux_inst_473: MUX2
        port map (
            O => mux_o_473,
            I0 => mux_o_437,
            I1 => mux_o_438,
            S0 => ad(5)
        );

    mux_inst_474: MUX2
        port map (
            O => mux_o_474,
            I0 => mux_o_439,
            I1 => mux_o_440,
            S0 => ad(5)
        );

    mux_inst_475: MUX2
        port map (
            O => mux_o_475,
            I0 => mux_o_441,
            I1 => mux_o_442,
            S0 => ad(5)
        );

    mux_inst_476: MUX2
        port map (
            O => mux_o_476,
            I0 => mux_o_443,
            I1 => mux_o_444,
            S0 => ad(5)
        );

    mux_inst_477: MUX2
        port map (
            O => mux_o_477,
            I0 => mux_o_445,
            I1 => mux_o_446,
            S0 => ad(6)
        );

    mux_inst_478: MUX2
        port map (
            O => mux_o_478,
            I0 => mux_o_447,
            I1 => mux_o_448,
            S0 => ad(6)
        );

    mux_inst_479: MUX2
        port map (
            O => mux_o_479,
            I0 => mux_o_449,
            I1 => mux_o_450,
            S0 => ad(6)
        );

    mux_inst_480: MUX2
        port map (
            O => mux_o_480,
            I0 => mux_o_451,
            I1 => mux_o_452,
            S0 => ad(6)
        );

    mux_inst_481: MUX2
        port map (
            O => mux_o_481,
            I0 => mux_o_453,
            I1 => mux_o_454,
            S0 => ad(6)
        );

    mux_inst_482: MUX2
        port map (
            O => mux_o_482,
            I0 => mux_o_455,
            I1 => mux_o_456,
            S0 => ad(6)
        );

    mux_inst_483: MUX2
        port map (
            O => mux_o_483,
            I0 => mux_o_457,
            I1 => mux_o_458,
            S0 => ad(6)
        );

    mux_inst_484: MUX2
        port map (
            O => mux_o_484,
            I0 => mux_o_459,
            I1 => mux_o_460,
            S0 => ad(6)
        );

    mux_inst_485: MUX2
        port map (
            O => mux_o_485,
            I0 => mux_o_461,
            I1 => mux_o_462,
            S0 => ad(6)
        );

    mux_inst_486: MUX2
        port map (
            O => mux_o_486,
            I0 => mux_o_463,
            I1 => mux_o_464,
            S0 => ad(6)
        );

    mux_inst_487: MUX2
        port map (
            O => mux_o_487,
            I0 => mux_o_465,
            I1 => mux_o_466,
            S0 => ad(6)
        );

    mux_inst_488: MUX2
        port map (
            O => mux_o_488,
            I0 => mux_o_467,
            I1 => mux_o_468,
            S0 => ad(6)
        );

    mux_inst_489: MUX2
        port map (
            O => mux_o_489,
            I0 => mux_o_469,
            I1 => mux_o_470,
            S0 => ad(6)
        );

    mux_inst_490: MUX2
        port map (
            O => mux_o_490,
            I0 => mux_o_471,
            I1 => mux_o_472,
            S0 => ad(6)
        );

    mux_inst_491: MUX2
        port map (
            O => mux_o_491,
            I0 => mux_o_473,
            I1 => mux_o_474,
            S0 => ad(6)
        );

    mux_inst_492: MUX2
        port map (
            O => mux_o_492,
            I0 => mux_o_475,
            I1 => mux_o_476,
            S0 => ad(6)
        );

    mux_inst_493: MUX2
        port map (
            O => mux_o_493,
            I0 => mux_o_477,
            I1 => mux_o_478,
            S0 => ad(7)
        );

    mux_inst_494: MUX2
        port map (
            O => mux_o_494,
            I0 => mux_o_479,
            I1 => mux_o_480,
            S0 => ad(7)
        );

    mux_inst_495: MUX2
        port map (
            O => mux_o_495,
            I0 => mux_o_481,
            I1 => mux_o_482,
            S0 => ad(7)
        );

    mux_inst_496: MUX2
        port map (
            O => mux_o_496,
            I0 => mux_o_483,
            I1 => mux_o_484,
            S0 => ad(7)
        );

    mux_inst_497: MUX2
        port map (
            O => mux_o_497,
            I0 => mux_o_485,
            I1 => mux_o_486,
            S0 => ad(7)
        );

    mux_inst_498: MUX2
        port map (
            O => mux_o_498,
            I0 => mux_o_487,
            I1 => mux_o_488,
            S0 => ad(7)
        );

    mux_inst_499: MUX2
        port map (
            O => mux_o_499,
            I0 => mux_o_489,
            I1 => mux_o_490,
            S0 => ad(7)
        );

    mux_inst_500: MUX2
        port map (
            O => mux_o_500,
            I0 => mux_o_491,
            I1 => mux_o_492,
            S0 => ad(7)
        );

    mux_inst_501: MUX2
        port map (
            O => mux_o_501,
            I0 => mux_o_493,
            I1 => mux_o_494,
            S0 => ad(8)
        );

    mux_inst_502: MUX2
        port map (
            O => mux_o_502,
            I0 => mux_o_495,
            I1 => mux_o_496,
            S0 => ad(8)
        );

    mux_inst_503: MUX2
        port map (
            O => mux_o_503,
            I0 => mux_o_497,
            I1 => mux_o_498,
            S0 => ad(8)
        );

    mux_inst_504: MUX2
        port map (
            O => mux_o_504,
            I0 => mux_o_499,
            I1 => mux_o_500,
            S0 => ad(8)
        );

    mux_inst_505: MUX2
        port map (
            O => mux_o_505,
            I0 => mux_o_501,
            I1 => mux_o_502,
            S0 => ad(9)
        );

    mux_inst_506: MUX2
        port map (
            O => mux_o_506,
            I0 => mux_o_503,
            I1 => mux_o_504,
            S0 => ad(9)
        );

    mux_inst_507: MUX2
        port map (
            O => dout(3),
            I0 => mux_o_505,
            I1 => mux_o_506,
            S0 => ad(10)
        );

    mux_inst_508: MUX2
        port map (
            O => mux_o_508,
            I0 => ram16s_inst_1_dout(4),
            I1 => ram16s_inst_3_dout(4),
            S0 => ad(4)
        );

    mux_inst_509: MUX2
        port map (
            O => mux_o_509,
            I0 => ram16s_inst_5_dout(4),
            I1 => ram16s_inst_7_dout(4),
            S0 => ad(4)
        );

    mux_inst_510: MUX2
        port map (
            O => mux_o_510,
            I0 => ram16s_inst_9_dout(4),
            I1 => ram16s_inst_11_dout(4),
            S0 => ad(4)
        );

    mux_inst_511: MUX2
        port map (
            O => mux_o_511,
            I0 => ram16s_inst_13_dout(4),
            I1 => ram16s_inst_15_dout(4),
            S0 => ad(4)
        );

    mux_inst_512: MUX2
        port map (
            O => mux_o_512,
            I0 => ram16s_inst_17_dout(4),
            I1 => ram16s_inst_19_dout(4),
            S0 => ad(4)
        );

    mux_inst_513: MUX2
        port map (
            O => mux_o_513,
            I0 => ram16s_inst_21_dout(4),
            I1 => ram16s_inst_23_dout(4),
            S0 => ad(4)
        );

    mux_inst_514: MUX2
        port map (
            O => mux_o_514,
            I0 => ram16s_inst_25_dout(4),
            I1 => ram16s_inst_27_dout(4),
            S0 => ad(4)
        );

    mux_inst_515: MUX2
        port map (
            O => mux_o_515,
            I0 => ram16s_inst_29_dout(4),
            I1 => ram16s_inst_31_dout(4),
            S0 => ad(4)
        );

    mux_inst_516: MUX2
        port map (
            O => mux_o_516,
            I0 => ram16s_inst_33_dout(4),
            I1 => ram16s_inst_35_dout(4),
            S0 => ad(4)
        );

    mux_inst_517: MUX2
        port map (
            O => mux_o_517,
            I0 => ram16s_inst_37_dout(4),
            I1 => ram16s_inst_39_dout(4),
            S0 => ad(4)
        );

    mux_inst_518: MUX2
        port map (
            O => mux_o_518,
            I0 => ram16s_inst_41_dout(4),
            I1 => ram16s_inst_43_dout(4),
            S0 => ad(4)
        );

    mux_inst_519: MUX2
        port map (
            O => mux_o_519,
            I0 => ram16s_inst_45_dout(4),
            I1 => ram16s_inst_47_dout(4),
            S0 => ad(4)
        );

    mux_inst_520: MUX2
        port map (
            O => mux_o_520,
            I0 => ram16s_inst_49_dout(4),
            I1 => ram16s_inst_51_dout(4),
            S0 => ad(4)
        );

    mux_inst_521: MUX2
        port map (
            O => mux_o_521,
            I0 => ram16s_inst_53_dout(4),
            I1 => ram16s_inst_55_dout(4),
            S0 => ad(4)
        );

    mux_inst_522: MUX2
        port map (
            O => mux_o_522,
            I0 => ram16s_inst_57_dout(4),
            I1 => ram16s_inst_59_dout(4),
            S0 => ad(4)
        );

    mux_inst_523: MUX2
        port map (
            O => mux_o_523,
            I0 => ram16s_inst_61_dout(4),
            I1 => ram16s_inst_63_dout(4),
            S0 => ad(4)
        );

    mux_inst_524: MUX2
        port map (
            O => mux_o_524,
            I0 => ram16s_inst_65_dout(4),
            I1 => ram16s_inst_67_dout(4),
            S0 => ad(4)
        );

    mux_inst_525: MUX2
        port map (
            O => mux_o_525,
            I0 => ram16s_inst_69_dout(4),
            I1 => ram16s_inst_71_dout(4),
            S0 => ad(4)
        );

    mux_inst_526: MUX2
        port map (
            O => mux_o_526,
            I0 => ram16s_inst_73_dout(4),
            I1 => ram16s_inst_75_dout(4),
            S0 => ad(4)
        );

    mux_inst_527: MUX2
        port map (
            O => mux_o_527,
            I0 => ram16s_inst_77_dout(4),
            I1 => ram16s_inst_79_dout(4),
            S0 => ad(4)
        );

    mux_inst_528: MUX2
        port map (
            O => mux_o_528,
            I0 => ram16s_inst_81_dout(4),
            I1 => ram16s_inst_83_dout(4),
            S0 => ad(4)
        );

    mux_inst_529: MUX2
        port map (
            O => mux_o_529,
            I0 => ram16s_inst_85_dout(4),
            I1 => ram16s_inst_87_dout(4),
            S0 => ad(4)
        );

    mux_inst_530: MUX2
        port map (
            O => mux_o_530,
            I0 => ram16s_inst_89_dout(4),
            I1 => ram16s_inst_91_dout(4),
            S0 => ad(4)
        );

    mux_inst_531: MUX2
        port map (
            O => mux_o_531,
            I0 => ram16s_inst_93_dout(4),
            I1 => ram16s_inst_95_dout(4),
            S0 => ad(4)
        );

    mux_inst_532: MUX2
        port map (
            O => mux_o_532,
            I0 => ram16s_inst_97_dout(4),
            I1 => ram16s_inst_99_dout(4),
            S0 => ad(4)
        );

    mux_inst_533: MUX2
        port map (
            O => mux_o_533,
            I0 => ram16s_inst_101_dout(4),
            I1 => ram16s_inst_103_dout(4),
            S0 => ad(4)
        );

    mux_inst_534: MUX2
        port map (
            O => mux_o_534,
            I0 => ram16s_inst_105_dout(4),
            I1 => ram16s_inst_107_dout(4),
            S0 => ad(4)
        );

    mux_inst_535: MUX2
        port map (
            O => mux_o_535,
            I0 => ram16s_inst_109_dout(4),
            I1 => ram16s_inst_111_dout(4),
            S0 => ad(4)
        );

    mux_inst_536: MUX2
        port map (
            O => mux_o_536,
            I0 => ram16s_inst_113_dout(4),
            I1 => ram16s_inst_115_dout(4),
            S0 => ad(4)
        );

    mux_inst_537: MUX2
        port map (
            O => mux_o_537,
            I0 => ram16s_inst_117_dout(4),
            I1 => ram16s_inst_119_dout(4),
            S0 => ad(4)
        );

    mux_inst_538: MUX2
        port map (
            O => mux_o_538,
            I0 => ram16s_inst_121_dout(4),
            I1 => ram16s_inst_123_dout(4),
            S0 => ad(4)
        );

    mux_inst_539: MUX2
        port map (
            O => mux_o_539,
            I0 => ram16s_inst_125_dout(4),
            I1 => ram16s_inst_127_dout(4),
            S0 => ad(4)
        );

    mux_inst_540: MUX2
        port map (
            O => mux_o_540,
            I0 => ram16s_inst_129_dout(4),
            I1 => ram16s_inst_131_dout(4),
            S0 => ad(4)
        );

    mux_inst_541: MUX2
        port map (
            O => mux_o_541,
            I0 => ram16s_inst_133_dout(4),
            I1 => ram16s_inst_135_dout(4),
            S0 => ad(4)
        );

    mux_inst_542: MUX2
        port map (
            O => mux_o_542,
            I0 => ram16s_inst_137_dout(4),
            I1 => ram16s_inst_139_dout(4),
            S0 => ad(4)
        );

    mux_inst_543: MUX2
        port map (
            O => mux_o_543,
            I0 => ram16s_inst_141_dout(4),
            I1 => ram16s_inst_143_dout(4),
            S0 => ad(4)
        );

    mux_inst_544: MUX2
        port map (
            O => mux_o_544,
            I0 => ram16s_inst_145_dout(4),
            I1 => ram16s_inst_147_dout(4),
            S0 => ad(4)
        );

    mux_inst_545: MUX2
        port map (
            O => mux_o_545,
            I0 => ram16s_inst_149_dout(4),
            I1 => ram16s_inst_151_dout(4),
            S0 => ad(4)
        );

    mux_inst_546: MUX2
        port map (
            O => mux_o_546,
            I0 => ram16s_inst_153_dout(4),
            I1 => ram16s_inst_155_dout(4),
            S0 => ad(4)
        );

    mux_inst_547: MUX2
        port map (
            O => mux_o_547,
            I0 => ram16s_inst_157_dout(4),
            I1 => ram16s_inst_159_dout(4),
            S0 => ad(4)
        );

    mux_inst_548: MUX2
        port map (
            O => mux_o_548,
            I0 => ram16s_inst_161_dout(4),
            I1 => ram16s_inst_163_dout(4),
            S0 => ad(4)
        );

    mux_inst_549: MUX2
        port map (
            O => mux_o_549,
            I0 => ram16s_inst_165_dout(4),
            I1 => ram16s_inst_167_dout(4),
            S0 => ad(4)
        );

    mux_inst_550: MUX2
        port map (
            O => mux_o_550,
            I0 => ram16s_inst_169_dout(4),
            I1 => ram16s_inst_171_dout(4),
            S0 => ad(4)
        );

    mux_inst_551: MUX2
        port map (
            O => mux_o_551,
            I0 => ram16s_inst_173_dout(4),
            I1 => ram16s_inst_175_dout(4),
            S0 => ad(4)
        );

    mux_inst_552: MUX2
        port map (
            O => mux_o_552,
            I0 => ram16s_inst_177_dout(4),
            I1 => ram16s_inst_179_dout(4),
            S0 => ad(4)
        );

    mux_inst_553: MUX2
        port map (
            O => mux_o_553,
            I0 => ram16s_inst_181_dout(4),
            I1 => ram16s_inst_183_dout(4),
            S0 => ad(4)
        );

    mux_inst_554: MUX2
        port map (
            O => mux_o_554,
            I0 => ram16s_inst_185_dout(4),
            I1 => ram16s_inst_187_dout(4),
            S0 => ad(4)
        );

    mux_inst_555: MUX2
        port map (
            O => mux_o_555,
            I0 => ram16s_inst_189_dout(4),
            I1 => ram16s_inst_191_dout(4),
            S0 => ad(4)
        );

    mux_inst_556: MUX2
        port map (
            O => mux_o_556,
            I0 => ram16s_inst_193_dout(4),
            I1 => ram16s_inst_195_dout(4),
            S0 => ad(4)
        );

    mux_inst_557: MUX2
        port map (
            O => mux_o_557,
            I0 => ram16s_inst_197_dout(4),
            I1 => ram16s_inst_199_dout(4),
            S0 => ad(4)
        );

    mux_inst_558: MUX2
        port map (
            O => mux_o_558,
            I0 => ram16s_inst_201_dout(4),
            I1 => ram16s_inst_203_dout(4),
            S0 => ad(4)
        );

    mux_inst_559: MUX2
        port map (
            O => mux_o_559,
            I0 => ram16s_inst_205_dout(4),
            I1 => ram16s_inst_207_dout(4),
            S0 => ad(4)
        );

    mux_inst_560: MUX2
        port map (
            O => mux_o_560,
            I0 => ram16s_inst_209_dout(4),
            I1 => ram16s_inst_211_dout(4),
            S0 => ad(4)
        );

    mux_inst_561: MUX2
        port map (
            O => mux_o_561,
            I0 => ram16s_inst_213_dout(4),
            I1 => ram16s_inst_215_dout(4),
            S0 => ad(4)
        );

    mux_inst_562: MUX2
        port map (
            O => mux_o_562,
            I0 => ram16s_inst_217_dout(4),
            I1 => ram16s_inst_219_dout(4),
            S0 => ad(4)
        );

    mux_inst_563: MUX2
        port map (
            O => mux_o_563,
            I0 => ram16s_inst_221_dout(4),
            I1 => ram16s_inst_223_dout(4),
            S0 => ad(4)
        );

    mux_inst_564: MUX2
        port map (
            O => mux_o_564,
            I0 => ram16s_inst_225_dout(4),
            I1 => ram16s_inst_227_dout(4),
            S0 => ad(4)
        );

    mux_inst_565: MUX2
        port map (
            O => mux_o_565,
            I0 => ram16s_inst_229_dout(4),
            I1 => ram16s_inst_231_dout(4),
            S0 => ad(4)
        );

    mux_inst_566: MUX2
        port map (
            O => mux_o_566,
            I0 => ram16s_inst_233_dout(4),
            I1 => ram16s_inst_235_dout(4),
            S0 => ad(4)
        );

    mux_inst_567: MUX2
        port map (
            O => mux_o_567,
            I0 => ram16s_inst_237_dout(4),
            I1 => ram16s_inst_239_dout(4),
            S0 => ad(4)
        );

    mux_inst_568: MUX2
        port map (
            O => mux_o_568,
            I0 => ram16s_inst_241_dout(4),
            I1 => ram16s_inst_243_dout(4),
            S0 => ad(4)
        );

    mux_inst_569: MUX2
        port map (
            O => mux_o_569,
            I0 => ram16s_inst_245_dout(4),
            I1 => ram16s_inst_247_dout(4),
            S0 => ad(4)
        );

    mux_inst_570: MUX2
        port map (
            O => mux_o_570,
            I0 => ram16s_inst_249_dout(4),
            I1 => ram16s_inst_251_dout(4),
            S0 => ad(4)
        );

    mux_inst_571: MUX2
        port map (
            O => mux_o_571,
            I0 => ram16s_inst_253_dout(4),
            I1 => ram16s_inst_255_dout(4),
            S0 => ad(4)
        );

    mux_inst_572: MUX2
        port map (
            O => mux_o_572,
            I0 => mux_o_508,
            I1 => mux_o_509,
            S0 => ad(5)
        );

    mux_inst_573: MUX2
        port map (
            O => mux_o_573,
            I0 => mux_o_510,
            I1 => mux_o_511,
            S0 => ad(5)
        );

    mux_inst_574: MUX2
        port map (
            O => mux_o_574,
            I0 => mux_o_512,
            I1 => mux_o_513,
            S0 => ad(5)
        );

    mux_inst_575: MUX2
        port map (
            O => mux_o_575,
            I0 => mux_o_514,
            I1 => mux_o_515,
            S0 => ad(5)
        );

    mux_inst_576: MUX2
        port map (
            O => mux_o_576,
            I0 => mux_o_516,
            I1 => mux_o_517,
            S0 => ad(5)
        );

    mux_inst_577: MUX2
        port map (
            O => mux_o_577,
            I0 => mux_o_518,
            I1 => mux_o_519,
            S0 => ad(5)
        );

    mux_inst_578: MUX2
        port map (
            O => mux_o_578,
            I0 => mux_o_520,
            I1 => mux_o_521,
            S0 => ad(5)
        );

    mux_inst_579: MUX2
        port map (
            O => mux_o_579,
            I0 => mux_o_522,
            I1 => mux_o_523,
            S0 => ad(5)
        );

    mux_inst_580: MUX2
        port map (
            O => mux_o_580,
            I0 => mux_o_524,
            I1 => mux_o_525,
            S0 => ad(5)
        );

    mux_inst_581: MUX2
        port map (
            O => mux_o_581,
            I0 => mux_o_526,
            I1 => mux_o_527,
            S0 => ad(5)
        );

    mux_inst_582: MUX2
        port map (
            O => mux_o_582,
            I0 => mux_o_528,
            I1 => mux_o_529,
            S0 => ad(5)
        );

    mux_inst_583: MUX2
        port map (
            O => mux_o_583,
            I0 => mux_o_530,
            I1 => mux_o_531,
            S0 => ad(5)
        );

    mux_inst_584: MUX2
        port map (
            O => mux_o_584,
            I0 => mux_o_532,
            I1 => mux_o_533,
            S0 => ad(5)
        );

    mux_inst_585: MUX2
        port map (
            O => mux_o_585,
            I0 => mux_o_534,
            I1 => mux_o_535,
            S0 => ad(5)
        );

    mux_inst_586: MUX2
        port map (
            O => mux_o_586,
            I0 => mux_o_536,
            I1 => mux_o_537,
            S0 => ad(5)
        );

    mux_inst_587: MUX2
        port map (
            O => mux_o_587,
            I0 => mux_o_538,
            I1 => mux_o_539,
            S0 => ad(5)
        );

    mux_inst_588: MUX2
        port map (
            O => mux_o_588,
            I0 => mux_o_540,
            I1 => mux_o_541,
            S0 => ad(5)
        );

    mux_inst_589: MUX2
        port map (
            O => mux_o_589,
            I0 => mux_o_542,
            I1 => mux_o_543,
            S0 => ad(5)
        );

    mux_inst_590: MUX2
        port map (
            O => mux_o_590,
            I0 => mux_o_544,
            I1 => mux_o_545,
            S0 => ad(5)
        );

    mux_inst_591: MUX2
        port map (
            O => mux_o_591,
            I0 => mux_o_546,
            I1 => mux_o_547,
            S0 => ad(5)
        );

    mux_inst_592: MUX2
        port map (
            O => mux_o_592,
            I0 => mux_o_548,
            I1 => mux_o_549,
            S0 => ad(5)
        );

    mux_inst_593: MUX2
        port map (
            O => mux_o_593,
            I0 => mux_o_550,
            I1 => mux_o_551,
            S0 => ad(5)
        );

    mux_inst_594: MUX2
        port map (
            O => mux_o_594,
            I0 => mux_o_552,
            I1 => mux_o_553,
            S0 => ad(5)
        );

    mux_inst_595: MUX2
        port map (
            O => mux_o_595,
            I0 => mux_o_554,
            I1 => mux_o_555,
            S0 => ad(5)
        );

    mux_inst_596: MUX2
        port map (
            O => mux_o_596,
            I0 => mux_o_556,
            I1 => mux_o_557,
            S0 => ad(5)
        );

    mux_inst_597: MUX2
        port map (
            O => mux_o_597,
            I0 => mux_o_558,
            I1 => mux_o_559,
            S0 => ad(5)
        );

    mux_inst_598: MUX2
        port map (
            O => mux_o_598,
            I0 => mux_o_560,
            I1 => mux_o_561,
            S0 => ad(5)
        );

    mux_inst_599: MUX2
        port map (
            O => mux_o_599,
            I0 => mux_o_562,
            I1 => mux_o_563,
            S0 => ad(5)
        );

    mux_inst_600: MUX2
        port map (
            O => mux_o_600,
            I0 => mux_o_564,
            I1 => mux_o_565,
            S0 => ad(5)
        );

    mux_inst_601: MUX2
        port map (
            O => mux_o_601,
            I0 => mux_o_566,
            I1 => mux_o_567,
            S0 => ad(5)
        );

    mux_inst_602: MUX2
        port map (
            O => mux_o_602,
            I0 => mux_o_568,
            I1 => mux_o_569,
            S0 => ad(5)
        );

    mux_inst_603: MUX2
        port map (
            O => mux_o_603,
            I0 => mux_o_570,
            I1 => mux_o_571,
            S0 => ad(5)
        );

    mux_inst_604: MUX2
        port map (
            O => mux_o_604,
            I0 => mux_o_572,
            I1 => mux_o_573,
            S0 => ad(6)
        );

    mux_inst_605: MUX2
        port map (
            O => mux_o_605,
            I0 => mux_o_574,
            I1 => mux_o_575,
            S0 => ad(6)
        );

    mux_inst_606: MUX2
        port map (
            O => mux_o_606,
            I0 => mux_o_576,
            I1 => mux_o_577,
            S0 => ad(6)
        );

    mux_inst_607: MUX2
        port map (
            O => mux_o_607,
            I0 => mux_o_578,
            I1 => mux_o_579,
            S0 => ad(6)
        );

    mux_inst_608: MUX2
        port map (
            O => mux_o_608,
            I0 => mux_o_580,
            I1 => mux_o_581,
            S0 => ad(6)
        );

    mux_inst_609: MUX2
        port map (
            O => mux_o_609,
            I0 => mux_o_582,
            I1 => mux_o_583,
            S0 => ad(6)
        );

    mux_inst_610: MUX2
        port map (
            O => mux_o_610,
            I0 => mux_o_584,
            I1 => mux_o_585,
            S0 => ad(6)
        );

    mux_inst_611: MUX2
        port map (
            O => mux_o_611,
            I0 => mux_o_586,
            I1 => mux_o_587,
            S0 => ad(6)
        );

    mux_inst_612: MUX2
        port map (
            O => mux_o_612,
            I0 => mux_o_588,
            I1 => mux_o_589,
            S0 => ad(6)
        );

    mux_inst_613: MUX2
        port map (
            O => mux_o_613,
            I0 => mux_o_590,
            I1 => mux_o_591,
            S0 => ad(6)
        );

    mux_inst_614: MUX2
        port map (
            O => mux_o_614,
            I0 => mux_o_592,
            I1 => mux_o_593,
            S0 => ad(6)
        );

    mux_inst_615: MUX2
        port map (
            O => mux_o_615,
            I0 => mux_o_594,
            I1 => mux_o_595,
            S0 => ad(6)
        );

    mux_inst_616: MUX2
        port map (
            O => mux_o_616,
            I0 => mux_o_596,
            I1 => mux_o_597,
            S0 => ad(6)
        );

    mux_inst_617: MUX2
        port map (
            O => mux_o_617,
            I0 => mux_o_598,
            I1 => mux_o_599,
            S0 => ad(6)
        );

    mux_inst_618: MUX2
        port map (
            O => mux_o_618,
            I0 => mux_o_600,
            I1 => mux_o_601,
            S0 => ad(6)
        );

    mux_inst_619: MUX2
        port map (
            O => mux_o_619,
            I0 => mux_o_602,
            I1 => mux_o_603,
            S0 => ad(6)
        );

    mux_inst_620: MUX2
        port map (
            O => mux_o_620,
            I0 => mux_o_604,
            I1 => mux_o_605,
            S0 => ad(7)
        );

    mux_inst_621: MUX2
        port map (
            O => mux_o_621,
            I0 => mux_o_606,
            I1 => mux_o_607,
            S0 => ad(7)
        );

    mux_inst_622: MUX2
        port map (
            O => mux_o_622,
            I0 => mux_o_608,
            I1 => mux_o_609,
            S0 => ad(7)
        );

    mux_inst_623: MUX2
        port map (
            O => mux_o_623,
            I0 => mux_o_610,
            I1 => mux_o_611,
            S0 => ad(7)
        );

    mux_inst_624: MUX2
        port map (
            O => mux_o_624,
            I0 => mux_o_612,
            I1 => mux_o_613,
            S0 => ad(7)
        );

    mux_inst_625: MUX2
        port map (
            O => mux_o_625,
            I0 => mux_o_614,
            I1 => mux_o_615,
            S0 => ad(7)
        );

    mux_inst_626: MUX2
        port map (
            O => mux_o_626,
            I0 => mux_o_616,
            I1 => mux_o_617,
            S0 => ad(7)
        );

    mux_inst_627: MUX2
        port map (
            O => mux_o_627,
            I0 => mux_o_618,
            I1 => mux_o_619,
            S0 => ad(7)
        );

    mux_inst_628: MUX2
        port map (
            O => mux_o_628,
            I0 => mux_o_620,
            I1 => mux_o_621,
            S0 => ad(8)
        );

    mux_inst_629: MUX2
        port map (
            O => mux_o_629,
            I0 => mux_o_622,
            I1 => mux_o_623,
            S0 => ad(8)
        );

    mux_inst_630: MUX2
        port map (
            O => mux_o_630,
            I0 => mux_o_624,
            I1 => mux_o_625,
            S0 => ad(8)
        );

    mux_inst_631: MUX2
        port map (
            O => mux_o_631,
            I0 => mux_o_626,
            I1 => mux_o_627,
            S0 => ad(8)
        );

    mux_inst_632: MUX2
        port map (
            O => mux_o_632,
            I0 => mux_o_628,
            I1 => mux_o_629,
            S0 => ad(9)
        );

    mux_inst_633: MUX2
        port map (
            O => mux_o_633,
            I0 => mux_o_630,
            I1 => mux_o_631,
            S0 => ad(9)
        );

    mux_inst_634: MUX2
        port map (
            O => dout(4),
            I0 => mux_o_632,
            I1 => mux_o_633,
            S0 => ad(10)
        );

    mux_inst_635: MUX2
        port map (
            O => mux_o_635,
            I0 => ram16s_inst_1_dout(5),
            I1 => ram16s_inst_3_dout(5),
            S0 => ad(4)
        );

    mux_inst_636: MUX2
        port map (
            O => mux_o_636,
            I0 => ram16s_inst_5_dout(5),
            I1 => ram16s_inst_7_dout(5),
            S0 => ad(4)
        );

    mux_inst_637: MUX2
        port map (
            O => mux_o_637,
            I0 => ram16s_inst_9_dout(5),
            I1 => ram16s_inst_11_dout(5),
            S0 => ad(4)
        );

    mux_inst_638: MUX2
        port map (
            O => mux_o_638,
            I0 => ram16s_inst_13_dout(5),
            I1 => ram16s_inst_15_dout(5),
            S0 => ad(4)
        );

    mux_inst_639: MUX2
        port map (
            O => mux_o_639,
            I0 => ram16s_inst_17_dout(5),
            I1 => ram16s_inst_19_dout(5),
            S0 => ad(4)
        );

    mux_inst_640: MUX2
        port map (
            O => mux_o_640,
            I0 => ram16s_inst_21_dout(5),
            I1 => ram16s_inst_23_dout(5),
            S0 => ad(4)
        );

    mux_inst_641: MUX2
        port map (
            O => mux_o_641,
            I0 => ram16s_inst_25_dout(5),
            I1 => ram16s_inst_27_dout(5),
            S0 => ad(4)
        );

    mux_inst_642: MUX2
        port map (
            O => mux_o_642,
            I0 => ram16s_inst_29_dout(5),
            I1 => ram16s_inst_31_dout(5),
            S0 => ad(4)
        );

    mux_inst_643: MUX2
        port map (
            O => mux_o_643,
            I0 => ram16s_inst_33_dout(5),
            I1 => ram16s_inst_35_dout(5),
            S0 => ad(4)
        );

    mux_inst_644: MUX2
        port map (
            O => mux_o_644,
            I0 => ram16s_inst_37_dout(5),
            I1 => ram16s_inst_39_dout(5),
            S0 => ad(4)
        );

    mux_inst_645: MUX2
        port map (
            O => mux_o_645,
            I0 => ram16s_inst_41_dout(5),
            I1 => ram16s_inst_43_dout(5),
            S0 => ad(4)
        );

    mux_inst_646: MUX2
        port map (
            O => mux_o_646,
            I0 => ram16s_inst_45_dout(5),
            I1 => ram16s_inst_47_dout(5),
            S0 => ad(4)
        );

    mux_inst_647: MUX2
        port map (
            O => mux_o_647,
            I0 => ram16s_inst_49_dout(5),
            I1 => ram16s_inst_51_dout(5),
            S0 => ad(4)
        );

    mux_inst_648: MUX2
        port map (
            O => mux_o_648,
            I0 => ram16s_inst_53_dout(5),
            I1 => ram16s_inst_55_dout(5),
            S0 => ad(4)
        );

    mux_inst_649: MUX2
        port map (
            O => mux_o_649,
            I0 => ram16s_inst_57_dout(5),
            I1 => ram16s_inst_59_dout(5),
            S0 => ad(4)
        );

    mux_inst_650: MUX2
        port map (
            O => mux_o_650,
            I0 => ram16s_inst_61_dout(5),
            I1 => ram16s_inst_63_dout(5),
            S0 => ad(4)
        );

    mux_inst_651: MUX2
        port map (
            O => mux_o_651,
            I0 => ram16s_inst_65_dout(5),
            I1 => ram16s_inst_67_dout(5),
            S0 => ad(4)
        );

    mux_inst_652: MUX2
        port map (
            O => mux_o_652,
            I0 => ram16s_inst_69_dout(5),
            I1 => ram16s_inst_71_dout(5),
            S0 => ad(4)
        );

    mux_inst_653: MUX2
        port map (
            O => mux_o_653,
            I0 => ram16s_inst_73_dout(5),
            I1 => ram16s_inst_75_dout(5),
            S0 => ad(4)
        );

    mux_inst_654: MUX2
        port map (
            O => mux_o_654,
            I0 => ram16s_inst_77_dout(5),
            I1 => ram16s_inst_79_dout(5),
            S0 => ad(4)
        );

    mux_inst_655: MUX2
        port map (
            O => mux_o_655,
            I0 => ram16s_inst_81_dout(5),
            I1 => ram16s_inst_83_dout(5),
            S0 => ad(4)
        );

    mux_inst_656: MUX2
        port map (
            O => mux_o_656,
            I0 => ram16s_inst_85_dout(5),
            I1 => ram16s_inst_87_dout(5),
            S0 => ad(4)
        );

    mux_inst_657: MUX2
        port map (
            O => mux_o_657,
            I0 => ram16s_inst_89_dout(5),
            I1 => ram16s_inst_91_dout(5),
            S0 => ad(4)
        );

    mux_inst_658: MUX2
        port map (
            O => mux_o_658,
            I0 => ram16s_inst_93_dout(5),
            I1 => ram16s_inst_95_dout(5),
            S0 => ad(4)
        );

    mux_inst_659: MUX2
        port map (
            O => mux_o_659,
            I0 => ram16s_inst_97_dout(5),
            I1 => ram16s_inst_99_dout(5),
            S0 => ad(4)
        );

    mux_inst_660: MUX2
        port map (
            O => mux_o_660,
            I0 => ram16s_inst_101_dout(5),
            I1 => ram16s_inst_103_dout(5),
            S0 => ad(4)
        );

    mux_inst_661: MUX2
        port map (
            O => mux_o_661,
            I0 => ram16s_inst_105_dout(5),
            I1 => ram16s_inst_107_dout(5),
            S0 => ad(4)
        );

    mux_inst_662: MUX2
        port map (
            O => mux_o_662,
            I0 => ram16s_inst_109_dout(5),
            I1 => ram16s_inst_111_dout(5),
            S0 => ad(4)
        );

    mux_inst_663: MUX2
        port map (
            O => mux_o_663,
            I0 => ram16s_inst_113_dout(5),
            I1 => ram16s_inst_115_dout(5),
            S0 => ad(4)
        );

    mux_inst_664: MUX2
        port map (
            O => mux_o_664,
            I0 => ram16s_inst_117_dout(5),
            I1 => ram16s_inst_119_dout(5),
            S0 => ad(4)
        );

    mux_inst_665: MUX2
        port map (
            O => mux_o_665,
            I0 => ram16s_inst_121_dout(5),
            I1 => ram16s_inst_123_dout(5),
            S0 => ad(4)
        );

    mux_inst_666: MUX2
        port map (
            O => mux_o_666,
            I0 => ram16s_inst_125_dout(5),
            I1 => ram16s_inst_127_dout(5),
            S0 => ad(4)
        );

    mux_inst_667: MUX2
        port map (
            O => mux_o_667,
            I0 => ram16s_inst_129_dout(5),
            I1 => ram16s_inst_131_dout(5),
            S0 => ad(4)
        );

    mux_inst_668: MUX2
        port map (
            O => mux_o_668,
            I0 => ram16s_inst_133_dout(5),
            I1 => ram16s_inst_135_dout(5),
            S0 => ad(4)
        );

    mux_inst_669: MUX2
        port map (
            O => mux_o_669,
            I0 => ram16s_inst_137_dout(5),
            I1 => ram16s_inst_139_dout(5),
            S0 => ad(4)
        );

    mux_inst_670: MUX2
        port map (
            O => mux_o_670,
            I0 => ram16s_inst_141_dout(5),
            I1 => ram16s_inst_143_dout(5),
            S0 => ad(4)
        );

    mux_inst_671: MUX2
        port map (
            O => mux_o_671,
            I0 => ram16s_inst_145_dout(5),
            I1 => ram16s_inst_147_dout(5),
            S0 => ad(4)
        );

    mux_inst_672: MUX2
        port map (
            O => mux_o_672,
            I0 => ram16s_inst_149_dout(5),
            I1 => ram16s_inst_151_dout(5),
            S0 => ad(4)
        );

    mux_inst_673: MUX2
        port map (
            O => mux_o_673,
            I0 => ram16s_inst_153_dout(5),
            I1 => ram16s_inst_155_dout(5),
            S0 => ad(4)
        );

    mux_inst_674: MUX2
        port map (
            O => mux_o_674,
            I0 => ram16s_inst_157_dout(5),
            I1 => ram16s_inst_159_dout(5),
            S0 => ad(4)
        );

    mux_inst_675: MUX2
        port map (
            O => mux_o_675,
            I0 => ram16s_inst_161_dout(5),
            I1 => ram16s_inst_163_dout(5),
            S0 => ad(4)
        );

    mux_inst_676: MUX2
        port map (
            O => mux_o_676,
            I0 => ram16s_inst_165_dout(5),
            I1 => ram16s_inst_167_dout(5),
            S0 => ad(4)
        );

    mux_inst_677: MUX2
        port map (
            O => mux_o_677,
            I0 => ram16s_inst_169_dout(5),
            I1 => ram16s_inst_171_dout(5),
            S0 => ad(4)
        );

    mux_inst_678: MUX2
        port map (
            O => mux_o_678,
            I0 => ram16s_inst_173_dout(5),
            I1 => ram16s_inst_175_dout(5),
            S0 => ad(4)
        );

    mux_inst_679: MUX2
        port map (
            O => mux_o_679,
            I0 => ram16s_inst_177_dout(5),
            I1 => ram16s_inst_179_dout(5),
            S0 => ad(4)
        );

    mux_inst_680: MUX2
        port map (
            O => mux_o_680,
            I0 => ram16s_inst_181_dout(5),
            I1 => ram16s_inst_183_dout(5),
            S0 => ad(4)
        );

    mux_inst_681: MUX2
        port map (
            O => mux_o_681,
            I0 => ram16s_inst_185_dout(5),
            I1 => ram16s_inst_187_dout(5),
            S0 => ad(4)
        );

    mux_inst_682: MUX2
        port map (
            O => mux_o_682,
            I0 => ram16s_inst_189_dout(5),
            I1 => ram16s_inst_191_dout(5),
            S0 => ad(4)
        );

    mux_inst_683: MUX2
        port map (
            O => mux_o_683,
            I0 => ram16s_inst_193_dout(5),
            I1 => ram16s_inst_195_dout(5),
            S0 => ad(4)
        );

    mux_inst_684: MUX2
        port map (
            O => mux_o_684,
            I0 => ram16s_inst_197_dout(5),
            I1 => ram16s_inst_199_dout(5),
            S0 => ad(4)
        );

    mux_inst_685: MUX2
        port map (
            O => mux_o_685,
            I0 => ram16s_inst_201_dout(5),
            I1 => ram16s_inst_203_dout(5),
            S0 => ad(4)
        );

    mux_inst_686: MUX2
        port map (
            O => mux_o_686,
            I0 => ram16s_inst_205_dout(5),
            I1 => ram16s_inst_207_dout(5),
            S0 => ad(4)
        );

    mux_inst_687: MUX2
        port map (
            O => mux_o_687,
            I0 => ram16s_inst_209_dout(5),
            I1 => ram16s_inst_211_dout(5),
            S0 => ad(4)
        );

    mux_inst_688: MUX2
        port map (
            O => mux_o_688,
            I0 => ram16s_inst_213_dout(5),
            I1 => ram16s_inst_215_dout(5),
            S0 => ad(4)
        );

    mux_inst_689: MUX2
        port map (
            O => mux_o_689,
            I0 => ram16s_inst_217_dout(5),
            I1 => ram16s_inst_219_dout(5),
            S0 => ad(4)
        );

    mux_inst_690: MUX2
        port map (
            O => mux_o_690,
            I0 => ram16s_inst_221_dout(5),
            I1 => ram16s_inst_223_dout(5),
            S0 => ad(4)
        );

    mux_inst_691: MUX2
        port map (
            O => mux_o_691,
            I0 => ram16s_inst_225_dout(5),
            I1 => ram16s_inst_227_dout(5),
            S0 => ad(4)
        );

    mux_inst_692: MUX2
        port map (
            O => mux_o_692,
            I0 => ram16s_inst_229_dout(5),
            I1 => ram16s_inst_231_dout(5),
            S0 => ad(4)
        );

    mux_inst_693: MUX2
        port map (
            O => mux_o_693,
            I0 => ram16s_inst_233_dout(5),
            I1 => ram16s_inst_235_dout(5),
            S0 => ad(4)
        );

    mux_inst_694: MUX2
        port map (
            O => mux_o_694,
            I0 => ram16s_inst_237_dout(5),
            I1 => ram16s_inst_239_dout(5),
            S0 => ad(4)
        );

    mux_inst_695: MUX2
        port map (
            O => mux_o_695,
            I0 => ram16s_inst_241_dout(5),
            I1 => ram16s_inst_243_dout(5),
            S0 => ad(4)
        );

    mux_inst_696: MUX2
        port map (
            O => mux_o_696,
            I0 => ram16s_inst_245_dout(5),
            I1 => ram16s_inst_247_dout(5),
            S0 => ad(4)
        );

    mux_inst_697: MUX2
        port map (
            O => mux_o_697,
            I0 => ram16s_inst_249_dout(5),
            I1 => ram16s_inst_251_dout(5),
            S0 => ad(4)
        );

    mux_inst_698: MUX2
        port map (
            O => mux_o_698,
            I0 => ram16s_inst_253_dout(5),
            I1 => ram16s_inst_255_dout(5),
            S0 => ad(4)
        );

    mux_inst_699: MUX2
        port map (
            O => mux_o_699,
            I0 => mux_o_635,
            I1 => mux_o_636,
            S0 => ad(5)
        );

    mux_inst_700: MUX2
        port map (
            O => mux_o_700,
            I0 => mux_o_637,
            I1 => mux_o_638,
            S0 => ad(5)
        );

    mux_inst_701: MUX2
        port map (
            O => mux_o_701,
            I0 => mux_o_639,
            I1 => mux_o_640,
            S0 => ad(5)
        );

    mux_inst_702: MUX2
        port map (
            O => mux_o_702,
            I0 => mux_o_641,
            I1 => mux_o_642,
            S0 => ad(5)
        );

    mux_inst_703: MUX2
        port map (
            O => mux_o_703,
            I0 => mux_o_643,
            I1 => mux_o_644,
            S0 => ad(5)
        );

    mux_inst_704: MUX2
        port map (
            O => mux_o_704,
            I0 => mux_o_645,
            I1 => mux_o_646,
            S0 => ad(5)
        );

    mux_inst_705: MUX2
        port map (
            O => mux_o_705,
            I0 => mux_o_647,
            I1 => mux_o_648,
            S0 => ad(5)
        );

    mux_inst_706: MUX2
        port map (
            O => mux_o_706,
            I0 => mux_o_649,
            I1 => mux_o_650,
            S0 => ad(5)
        );

    mux_inst_707: MUX2
        port map (
            O => mux_o_707,
            I0 => mux_o_651,
            I1 => mux_o_652,
            S0 => ad(5)
        );

    mux_inst_708: MUX2
        port map (
            O => mux_o_708,
            I0 => mux_o_653,
            I1 => mux_o_654,
            S0 => ad(5)
        );

    mux_inst_709: MUX2
        port map (
            O => mux_o_709,
            I0 => mux_o_655,
            I1 => mux_o_656,
            S0 => ad(5)
        );

    mux_inst_710: MUX2
        port map (
            O => mux_o_710,
            I0 => mux_o_657,
            I1 => mux_o_658,
            S0 => ad(5)
        );

    mux_inst_711: MUX2
        port map (
            O => mux_o_711,
            I0 => mux_o_659,
            I1 => mux_o_660,
            S0 => ad(5)
        );

    mux_inst_712: MUX2
        port map (
            O => mux_o_712,
            I0 => mux_o_661,
            I1 => mux_o_662,
            S0 => ad(5)
        );

    mux_inst_713: MUX2
        port map (
            O => mux_o_713,
            I0 => mux_o_663,
            I1 => mux_o_664,
            S0 => ad(5)
        );

    mux_inst_714: MUX2
        port map (
            O => mux_o_714,
            I0 => mux_o_665,
            I1 => mux_o_666,
            S0 => ad(5)
        );

    mux_inst_715: MUX2
        port map (
            O => mux_o_715,
            I0 => mux_o_667,
            I1 => mux_o_668,
            S0 => ad(5)
        );

    mux_inst_716: MUX2
        port map (
            O => mux_o_716,
            I0 => mux_o_669,
            I1 => mux_o_670,
            S0 => ad(5)
        );

    mux_inst_717: MUX2
        port map (
            O => mux_o_717,
            I0 => mux_o_671,
            I1 => mux_o_672,
            S0 => ad(5)
        );

    mux_inst_718: MUX2
        port map (
            O => mux_o_718,
            I0 => mux_o_673,
            I1 => mux_o_674,
            S0 => ad(5)
        );

    mux_inst_719: MUX2
        port map (
            O => mux_o_719,
            I0 => mux_o_675,
            I1 => mux_o_676,
            S0 => ad(5)
        );

    mux_inst_720: MUX2
        port map (
            O => mux_o_720,
            I0 => mux_o_677,
            I1 => mux_o_678,
            S0 => ad(5)
        );

    mux_inst_721: MUX2
        port map (
            O => mux_o_721,
            I0 => mux_o_679,
            I1 => mux_o_680,
            S0 => ad(5)
        );

    mux_inst_722: MUX2
        port map (
            O => mux_o_722,
            I0 => mux_o_681,
            I1 => mux_o_682,
            S0 => ad(5)
        );

    mux_inst_723: MUX2
        port map (
            O => mux_o_723,
            I0 => mux_o_683,
            I1 => mux_o_684,
            S0 => ad(5)
        );

    mux_inst_724: MUX2
        port map (
            O => mux_o_724,
            I0 => mux_o_685,
            I1 => mux_o_686,
            S0 => ad(5)
        );

    mux_inst_725: MUX2
        port map (
            O => mux_o_725,
            I0 => mux_o_687,
            I1 => mux_o_688,
            S0 => ad(5)
        );

    mux_inst_726: MUX2
        port map (
            O => mux_o_726,
            I0 => mux_o_689,
            I1 => mux_o_690,
            S0 => ad(5)
        );

    mux_inst_727: MUX2
        port map (
            O => mux_o_727,
            I0 => mux_o_691,
            I1 => mux_o_692,
            S0 => ad(5)
        );

    mux_inst_728: MUX2
        port map (
            O => mux_o_728,
            I0 => mux_o_693,
            I1 => mux_o_694,
            S0 => ad(5)
        );

    mux_inst_729: MUX2
        port map (
            O => mux_o_729,
            I0 => mux_o_695,
            I1 => mux_o_696,
            S0 => ad(5)
        );

    mux_inst_730: MUX2
        port map (
            O => mux_o_730,
            I0 => mux_o_697,
            I1 => mux_o_698,
            S0 => ad(5)
        );

    mux_inst_731: MUX2
        port map (
            O => mux_o_731,
            I0 => mux_o_699,
            I1 => mux_o_700,
            S0 => ad(6)
        );

    mux_inst_732: MUX2
        port map (
            O => mux_o_732,
            I0 => mux_o_701,
            I1 => mux_o_702,
            S0 => ad(6)
        );

    mux_inst_733: MUX2
        port map (
            O => mux_o_733,
            I0 => mux_o_703,
            I1 => mux_o_704,
            S0 => ad(6)
        );

    mux_inst_734: MUX2
        port map (
            O => mux_o_734,
            I0 => mux_o_705,
            I1 => mux_o_706,
            S0 => ad(6)
        );

    mux_inst_735: MUX2
        port map (
            O => mux_o_735,
            I0 => mux_o_707,
            I1 => mux_o_708,
            S0 => ad(6)
        );

    mux_inst_736: MUX2
        port map (
            O => mux_o_736,
            I0 => mux_o_709,
            I1 => mux_o_710,
            S0 => ad(6)
        );

    mux_inst_737: MUX2
        port map (
            O => mux_o_737,
            I0 => mux_o_711,
            I1 => mux_o_712,
            S0 => ad(6)
        );

    mux_inst_738: MUX2
        port map (
            O => mux_o_738,
            I0 => mux_o_713,
            I1 => mux_o_714,
            S0 => ad(6)
        );

    mux_inst_739: MUX2
        port map (
            O => mux_o_739,
            I0 => mux_o_715,
            I1 => mux_o_716,
            S0 => ad(6)
        );

    mux_inst_740: MUX2
        port map (
            O => mux_o_740,
            I0 => mux_o_717,
            I1 => mux_o_718,
            S0 => ad(6)
        );

    mux_inst_741: MUX2
        port map (
            O => mux_o_741,
            I0 => mux_o_719,
            I1 => mux_o_720,
            S0 => ad(6)
        );

    mux_inst_742: MUX2
        port map (
            O => mux_o_742,
            I0 => mux_o_721,
            I1 => mux_o_722,
            S0 => ad(6)
        );

    mux_inst_743: MUX2
        port map (
            O => mux_o_743,
            I0 => mux_o_723,
            I1 => mux_o_724,
            S0 => ad(6)
        );

    mux_inst_744: MUX2
        port map (
            O => mux_o_744,
            I0 => mux_o_725,
            I1 => mux_o_726,
            S0 => ad(6)
        );

    mux_inst_745: MUX2
        port map (
            O => mux_o_745,
            I0 => mux_o_727,
            I1 => mux_o_728,
            S0 => ad(6)
        );

    mux_inst_746: MUX2
        port map (
            O => mux_o_746,
            I0 => mux_o_729,
            I1 => mux_o_730,
            S0 => ad(6)
        );

    mux_inst_747: MUX2
        port map (
            O => mux_o_747,
            I0 => mux_o_731,
            I1 => mux_o_732,
            S0 => ad(7)
        );

    mux_inst_748: MUX2
        port map (
            O => mux_o_748,
            I0 => mux_o_733,
            I1 => mux_o_734,
            S0 => ad(7)
        );

    mux_inst_749: MUX2
        port map (
            O => mux_o_749,
            I0 => mux_o_735,
            I1 => mux_o_736,
            S0 => ad(7)
        );

    mux_inst_750: MUX2
        port map (
            O => mux_o_750,
            I0 => mux_o_737,
            I1 => mux_o_738,
            S0 => ad(7)
        );

    mux_inst_751: MUX2
        port map (
            O => mux_o_751,
            I0 => mux_o_739,
            I1 => mux_o_740,
            S0 => ad(7)
        );

    mux_inst_752: MUX2
        port map (
            O => mux_o_752,
            I0 => mux_o_741,
            I1 => mux_o_742,
            S0 => ad(7)
        );

    mux_inst_753: MUX2
        port map (
            O => mux_o_753,
            I0 => mux_o_743,
            I1 => mux_o_744,
            S0 => ad(7)
        );

    mux_inst_754: MUX2
        port map (
            O => mux_o_754,
            I0 => mux_o_745,
            I1 => mux_o_746,
            S0 => ad(7)
        );

    mux_inst_755: MUX2
        port map (
            O => mux_o_755,
            I0 => mux_o_747,
            I1 => mux_o_748,
            S0 => ad(8)
        );

    mux_inst_756: MUX2
        port map (
            O => mux_o_756,
            I0 => mux_o_749,
            I1 => mux_o_750,
            S0 => ad(8)
        );

    mux_inst_757: MUX2
        port map (
            O => mux_o_757,
            I0 => mux_o_751,
            I1 => mux_o_752,
            S0 => ad(8)
        );

    mux_inst_758: MUX2
        port map (
            O => mux_o_758,
            I0 => mux_o_753,
            I1 => mux_o_754,
            S0 => ad(8)
        );

    mux_inst_759: MUX2
        port map (
            O => mux_o_759,
            I0 => mux_o_755,
            I1 => mux_o_756,
            S0 => ad(9)
        );

    mux_inst_760: MUX2
        port map (
            O => mux_o_760,
            I0 => mux_o_757,
            I1 => mux_o_758,
            S0 => ad(9)
        );

    mux_inst_761: MUX2
        port map (
            O => dout(5),
            I0 => mux_o_759,
            I1 => mux_o_760,
            S0 => ad(10)
        );

    mux_inst_762: MUX2
        port map (
            O => mux_o_762,
            I0 => ram16s_inst_1_dout(6),
            I1 => ram16s_inst_3_dout(6),
            S0 => ad(4)
        );

    mux_inst_763: MUX2
        port map (
            O => mux_o_763,
            I0 => ram16s_inst_5_dout(6),
            I1 => ram16s_inst_7_dout(6),
            S0 => ad(4)
        );

    mux_inst_764: MUX2
        port map (
            O => mux_o_764,
            I0 => ram16s_inst_9_dout(6),
            I1 => ram16s_inst_11_dout(6),
            S0 => ad(4)
        );

    mux_inst_765: MUX2
        port map (
            O => mux_o_765,
            I0 => ram16s_inst_13_dout(6),
            I1 => ram16s_inst_15_dout(6),
            S0 => ad(4)
        );

    mux_inst_766: MUX2
        port map (
            O => mux_o_766,
            I0 => ram16s_inst_17_dout(6),
            I1 => ram16s_inst_19_dout(6),
            S0 => ad(4)
        );

    mux_inst_767: MUX2
        port map (
            O => mux_o_767,
            I0 => ram16s_inst_21_dout(6),
            I1 => ram16s_inst_23_dout(6),
            S0 => ad(4)
        );

    mux_inst_768: MUX2
        port map (
            O => mux_o_768,
            I0 => ram16s_inst_25_dout(6),
            I1 => ram16s_inst_27_dout(6),
            S0 => ad(4)
        );

    mux_inst_769: MUX2
        port map (
            O => mux_o_769,
            I0 => ram16s_inst_29_dout(6),
            I1 => ram16s_inst_31_dout(6),
            S0 => ad(4)
        );

    mux_inst_770: MUX2
        port map (
            O => mux_o_770,
            I0 => ram16s_inst_33_dout(6),
            I1 => ram16s_inst_35_dout(6),
            S0 => ad(4)
        );

    mux_inst_771: MUX2
        port map (
            O => mux_o_771,
            I0 => ram16s_inst_37_dout(6),
            I1 => ram16s_inst_39_dout(6),
            S0 => ad(4)
        );

    mux_inst_772: MUX2
        port map (
            O => mux_o_772,
            I0 => ram16s_inst_41_dout(6),
            I1 => ram16s_inst_43_dout(6),
            S0 => ad(4)
        );

    mux_inst_773: MUX2
        port map (
            O => mux_o_773,
            I0 => ram16s_inst_45_dout(6),
            I1 => ram16s_inst_47_dout(6),
            S0 => ad(4)
        );

    mux_inst_774: MUX2
        port map (
            O => mux_o_774,
            I0 => ram16s_inst_49_dout(6),
            I1 => ram16s_inst_51_dout(6),
            S0 => ad(4)
        );

    mux_inst_775: MUX2
        port map (
            O => mux_o_775,
            I0 => ram16s_inst_53_dout(6),
            I1 => ram16s_inst_55_dout(6),
            S0 => ad(4)
        );

    mux_inst_776: MUX2
        port map (
            O => mux_o_776,
            I0 => ram16s_inst_57_dout(6),
            I1 => ram16s_inst_59_dout(6),
            S0 => ad(4)
        );

    mux_inst_777: MUX2
        port map (
            O => mux_o_777,
            I0 => ram16s_inst_61_dout(6),
            I1 => ram16s_inst_63_dout(6),
            S0 => ad(4)
        );

    mux_inst_778: MUX2
        port map (
            O => mux_o_778,
            I0 => ram16s_inst_65_dout(6),
            I1 => ram16s_inst_67_dout(6),
            S0 => ad(4)
        );

    mux_inst_779: MUX2
        port map (
            O => mux_o_779,
            I0 => ram16s_inst_69_dout(6),
            I1 => ram16s_inst_71_dout(6),
            S0 => ad(4)
        );

    mux_inst_780: MUX2
        port map (
            O => mux_o_780,
            I0 => ram16s_inst_73_dout(6),
            I1 => ram16s_inst_75_dout(6),
            S0 => ad(4)
        );

    mux_inst_781: MUX2
        port map (
            O => mux_o_781,
            I0 => ram16s_inst_77_dout(6),
            I1 => ram16s_inst_79_dout(6),
            S0 => ad(4)
        );

    mux_inst_782: MUX2
        port map (
            O => mux_o_782,
            I0 => ram16s_inst_81_dout(6),
            I1 => ram16s_inst_83_dout(6),
            S0 => ad(4)
        );

    mux_inst_783: MUX2
        port map (
            O => mux_o_783,
            I0 => ram16s_inst_85_dout(6),
            I1 => ram16s_inst_87_dout(6),
            S0 => ad(4)
        );

    mux_inst_784: MUX2
        port map (
            O => mux_o_784,
            I0 => ram16s_inst_89_dout(6),
            I1 => ram16s_inst_91_dout(6),
            S0 => ad(4)
        );

    mux_inst_785: MUX2
        port map (
            O => mux_o_785,
            I0 => ram16s_inst_93_dout(6),
            I1 => ram16s_inst_95_dout(6),
            S0 => ad(4)
        );

    mux_inst_786: MUX2
        port map (
            O => mux_o_786,
            I0 => ram16s_inst_97_dout(6),
            I1 => ram16s_inst_99_dout(6),
            S0 => ad(4)
        );

    mux_inst_787: MUX2
        port map (
            O => mux_o_787,
            I0 => ram16s_inst_101_dout(6),
            I1 => ram16s_inst_103_dout(6),
            S0 => ad(4)
        );

    mux_inst_788: MUX2
        port map (
            O => mux_o_788,
            I0 => ram16s_inst_105_dout(6),
            I1 => ram16s_inst_107_dout(6),
            S0 => ad(4)
        );

    mux_inst_789: MUX2
        port map (
            O => mux_o_789,
            I0 => ram16s_inst_109_dout(6),
            I1 => ram16s_inst_111_dout(6),
            S0 => ad(4)
        );

    mux_inst_790: MUX2
        port map (
            O => mux_o_790,
            I0 => ram16s_inst_113_dout(6),
            I1 => ram16s_inst_115_dout(6),
            S0 => ad(4)
        );

    mux_inst_791: MUX2
        port map (
            O => mux_o_791,
            I0 => ram16s_inst_117_dout(6),
            I1 => ram16s_inst_119_dout(6),
            S0 => ad(4)
        );

    mux_inst_792: MUX2
        port map (
            O => mux_o_792,
            I0 => ram16s_inst_121_dout(6),
            I1 => ram16s_inst_123_dout(6),
            S0 => ad(4)
        );

    mux_inst_793: MUX2
        port map (
            O => mux_o_793,
            I0 => ram16s_inst_125_dout(6),
            I1 => ram16s_inst_127_dout(6),
            S0 => ad(4)
        );

    mux_inst_794: MUX2
        port map (
            O => mux_o_794,
            I0 => ram16s_inst_129_dout(6),
            I1 => ram16s_inst_131_dout(6),
            S0 => ad(4)
        );

    mux_inst_795: MUX2
        port map (
            O => mux_o_795,
            I0 => ram16s_inst_133_dout(6),
            I1 => ram16s_inst_135_dout(6),
            S0 => ad(4)
        );

    mux_inst_796: MUX2
        port map (
            O => mux_o_796,
            I0 => ram16s_inst_137_dout(6),
            I1 => ram16s_inst_139_dout(6),
            S0 => ad(4)
        );

    mux_inst_797: MUX2
        port map (
            O => mux_o_797,
            I0 => ram16s_inst_141_dout(6),
            I1 => ram16s_inst_143_dout(6),
            S0 => ad(4)
        );

    mux_inst_798: MUX2
        port map (
            O => mux_o_798,
            I0 => ram16s_inst_145_dout(6),
            I1 => ram16s_inst_147_dout(6),
            S0 => ad(4)
        );

    mux_inst_799: MUX2
        port map (
            O => mux_o_799,
            I0 => ram16s_inst_149_dout(6),
            I1 => ram16s_inst_151_dout(6),
            S0 => ad(4)
        );

    mux_inst_800: MUX2
        port map (
            O => mux_o_800,
            I0 => ram16s_inst_153_dout(6),
            I1 => ram16s_inst_155_dout(6),
            S0 => ad(4)
        );

    mux_inst_801: MUX2
        port map (
            O => mux_o_801,
            I0 => ram16s_inst_157_dout(6),
            I1 => ram16s_inst_159_dout(6),
            S0 => ad(4)
        );

    mux_inst_802: MUX2
        port map (
            O => mux_o_802,
            I0 => ram16s_inst_161_dout(6),
            I1 => ram16s_inst_163_dout(6),
            S0 => ad(4)
        );

    mux_inst_803: MUX2
        port map (
            O => mux_o_803,
            I0 => ram16s_inst_165_dout(6),
            I1 => ram16s_inst_167_dout(6),
            S0 => ad(4)
        );

    mux_inst_804: MUX2
        port map (
            O => mux_o_804,
            I0 => ram16s_inst_169_dout(6),
            I1 => ram16s_inst_171_dout(6),
            S0 => ad(4)
        );

    mux_inst_805: MUX2
        port map (
            O => mux_o_805,
            I0 => ram16s_inst_173_dout(6),
            I1 => ram16s_inst_175_dout(6),
            S0 => ad(4)
        );

    mux_inst_806: MUX2
        port map (
            O => mux_o_806,
            I0 => ram16s_inst_177_dout(6),
            I1 => ram16s_inst_179_dout(6),
            S0 => ad(4)
        );

    mux_inst_807: MUX2
        port map (
            O => mux_o_807,
            I0 => ram16s_inst_181_dout(6),
            I1 => ram16s_inst_183_dout(6),
            S0 => ad(4)
        );

    mux_inst_808: MUX2
        port map (
            O => mux_o_808,
            I0 => ram16s_inst_185_dout(6),
            I1 => ram16s_inst_187_dout(6),
            S0 => ad(4)
        );

    mux_inst_809: MUX2
        port map (
            O => mux_o_809,
            I0 => ram16s_inst_189_dout(6),
            I1 => ram16s_inst_191_dout(6),
            S0 => ad(4)
        );

    mux_inst_810: MUX2
        port map (
            O => mux_o_810,
            I0 => ram16s_inst_193_dout(6),
            I1 => ram16s_inst_195_dout(6),
            S0 => ad(4)
        );

    mux_inst_811: MUX2
        port map (
            O => mux_o_811,
            I0 => ram16s_inst_197_dout(6),
            I1 => ram16s_inst_199_dout(6),
            S0 => ad(4)
        );

    mux_inst_812: MUX2
        port map (
            O => mux_o_812,
            I0 => ram16s_inst_201_dout(6),
            I1 => ram16s_inst_203_dout(6),
            S0 => ad(4)
        );

    mux_inst_813: MUX2
        port map (
            O => mux_o_813,
            I0 => ram16s_inst_205_dout(6),
            I1 => ram16s_inst_207_dout(6),
            S0 => ad(4)
        );

    mux_inst_814: MUX2
        port map (
            O => mux_o_814,
            I0 => ram16s_inst_209_dout(6),
            I1 => ram16s_inst_211_dout(6),
            S0 => ad(4)
        );

    mux_inst_815: MUX2
        port map (
            O => mux_o_815,
            I0 => ram16s_inst_213_dout(6),
            I1 => ram16s_inst_215_dout(6),
            S0 => ad(4)
        );

    mux_inst_816: MUX2
        port map (
            O => mux_o_816,
            I0 => ram16s_inst_217_dout(6),
            I1 => ram16s_inst_219_dout(6),
            S0 => ad(4)
        );

    mux_inst_817: MUX2
        port map (
            O => mux_o_817,
            I0 => ram16s_inst_221_dout(6),
            I1 => ram16s_inst_223_dout(6),
            S0 => ad(4)
        );

    mux_inst_818: MUX2
        port map (
            O => mux_o_818,
            I0 => ram16s_inst_225_dout(6),
            I1 => ram16s_inst_227_dout(6),
            S0 => ad(4)
        );

    mux_inst_819: MUX2
        port map (
            O => mux_o_819,
            I0 => ram16s_inst_229_dout(6),
            I1 => ram16s_inst_231_dout(6),
            S0 => ad(4)
        );

    mux_inst_820: MUX2
        port map (
            O => mux_o_820,
            I0 => ram16s_inst_233_dout(6),
            I1 => ram16s_inst_235_dout(6),
            S0 => ad(4)
        );

    mux_inst_821: MUX2
        port map (
            O => mux_o_821,
            I0 => ram16s_inst_237_dout(6),
            I1 => ram16s_inst_239_dout(6),
            S0 => ad(4)
        );

    mux_inst_822: MUX2
        port map (
            O => mux_o_822,
            I0 => ram16s_inst_241_dout(6),
            I1 => ram16s_inst_243_dout(6),
            S0 => ad(4)
        );

    mux_inst_823: MUX2
        port map (
            O => mux_o_823,
            I0 => ram16s_inst_245_dout(6),
            I1 => ram16s_inst_247_dout(6),
            S0 => ad(4)
        );

    mux_inst_824: MUX2
        port map (
            O => mux_o_824,
            I0 => ram16s_inst_249_dout(6),
            I1 => ram16s_inst_251_dout(6),
            S0 => ad(4)
        );

    mux_inst_825: MUX2
        port map (
            O => mux_o_825,
            I0 => ram16s_inst_253_dout(6),
            I1 => ram16s_inst_255_dout(6),
            S0 => ad(4)
        );

    mux_inst_826: MUX2
        port map (
            O => mux_o_826,
            I0 => mux_o_762,
            I1 => mux_o_763,
            S0 => ad(5)
        );

    mux_inst_827: MUX2
        port map (
            O => mux_o_827,
            I0 => mux_o_764,
            I1 => mux_o_765,
            S0 => ad(5)
        );

    mux_inst_828: MUX2
        port map (
            O => mux_o_828,
            I0 => mux_o_766,
            I1 => mux_o_767,
            S0 => ad(5)
        );

    mux_inst_829: MUX2
        port map (
            O => mux_o_829,
            I0 => mux_o_768,
            I1 => mux_o_769,
            S0 => ad(5)
        );

    mux_inst_830: MUX2
        port map (
            O => mux_o_830,
            I0 => mux_o_770,
            I1 => mux_o_771,
            S0 => ad(5)
        );

    mux_inst_831: MUX2
        port map (
            O => mux_o_831,
            I0 => mux_o_772,
            I1 => mux_o_773,
            S0 => ad(5)
        );

    mux_inst_832: MUX2
        port map (
            O => mux_o_832,
            I0 => mux_o_774,
            I1 => mux_o_775,
            S0 => ad(5)
        );

    mux_inst_833: MUX2
        port map (
            O => mux_o_833,
            I0 => mux_o_776,
            I1 => mux_o_777,
            S0 => ad(5)
        );

    mux_inst_834: MUX2
        port map (
            O => mux_o_834,
            I0 => mux_o_778,
            I1 => mux_o_779,
            S0 => ad(5)
        );

    mux_inst_835: MUX2
        port map (
            O => mux_o_835,
            I0 => mux_o_780,
            I1 => mux_o_781,
            S0 => ad(5)
        );

    mux_inst_836: MUX2
        port map (
            O => mux_o_836,
            I0 => mux_o_782,
            I1 => mux_o_783,
            S0 => ad(5)
        );

    mux_inst_837: MUX2
        port map (
            O => mux_o_837,
            I0 => mux_o_784,
            I1 => mux_o_785,
            S0 => ad(5)
        );

    mux_inst_838: MUX2
        port map (
            O => mux_o_838,
            I0 => mux_o_786,
            I1 => mux_o_787,
            S0 => ad(5)
        );

    mux_inst_839: MUX2
        port map (
            O => mux_o_839,
            I0 => mux_o_788,
            I1 => mux_o_789,
            S0 => ad(5)
        );

    mux_inst_840: MUX2
        port map (
            O => mux_o_840,
            I0 => mux_o_790,
            I1 => mux_o_791,
            S0 => ad(5)
        );

    mux_inst_841: MUX2
        port map (
            O => mux_o_841,
            I0 => mux_o_792,
            I1 => mux_o_793,
            S0 => ad(5)
        );

    mux_inst_842: MUX2
        port map (
            O => mux_o_842,
            I0 => mux_o_794,
            I1 => mux_o_795,
            S0 => ad(5)
        );

    mux_inst_843: MUX2
        port map (
            O => mux_o_843,
            I0 => mux_o_796,
            I1 => mux_o_797,
            S0 => ad(5)
        );

    mux_inst_844: MUX2
        port map (
            O => mux_o_844,
            I0 => mux_o_798,
            I1 => mux_o_799,
            S0 => ad(5)
        );

    mux_inst_845: MUX2
        port map (
            O => mux_o_845,
            I0 => mux_o_800,
            I1 => mux_o_801,
            S0 => ad(5)
        );

    mux_inst_846: MUX2
        port map (
            O => mux_o_846,
            I0 => mux_o_802,
            I1 => mux_o_803,
            S0 => ad(5)
        );

    mux_inst_847: MUX2
        port map (
            O => mux_o_847,
            I0 => mux_o_804,
            I1 => mux_o_805,
            S0 => ad(5)
        );

    mux_inst_848: MUX2
        port map (
            O => mux_o_848,
            I0 => mux_o_806,
            I1 => mux_o_807,
            S0 => ad(5)
        );

    mux_inst_849: MUX2
        port map (
            O => mux_o_849,
            I0 => mux_o_808,
            I1 => mux_o_809,
            S0 => ad(5)
        );

    mux_inst_850: MUX2
        port map (
            O => mux_o_850,
            I0 => mux_o_810,
            I1 => mux_o_811,
            S0 => ad(5)
        );

    mux_inst_851: MUX2
        port map (
            O => mux_o_851,
            I0 => mux_o_812,
            I1 => mux_o_813,
            S0 => ad(5)
        );

    mux_inst_852: MUX2
        port map (
            O => mux_o_852,
            I0 => mux_o_814,
            I1 => mux_o_815,
            S0 => ad(5)
        );

    mux_inst_853: MUX2
        port map (
            O => mux_o_853,
            I0 => mux_o_816,
            I1 => mux_o_817,
            S0 => ad(5)
        );

    mux_inst_854: MUX2
        port map (
            O => mux_o_854,
            I0 => mux_o_818,
            I1 => mux_o_819,
            S0 => ad(5)
        );

    mux_inst_855: MUX2
        port map (
            O => mux_o_855,
            I0 => mux_o_820,
            I1 => mux_o_821,
            S0 => ad(5)
        );

    mux_inst_856: MUX2
        port map (
            O => mux_o_856,
            I0 => mux_o_822,
            I1 => mux_o_823,
            S0 => ad(5)
        );

    mux_inst_857: MUX2
        port map (
            O => mux_o_857,
            I0 => mux_o_824,
            I1 => mux_o_825,
            S0 => ad(5)
        );

    mux_inst_858: MUX2
        port map (
            O => mux_o_858,
            I0 => mux_o_826,
            I1 => mux_o_827,
            S0 => ad(6)
        );

    mux_inst_859: MUX2
        port map (
            O => mux_o_859,
            I0 => mux_o_828,
            I1 => mux_o_829,
            S0 => ad(6)
        );

    mux_inst_860: MUX2
        port map (
            O => mux_o_860,
            I0 => mux_o_830,
            I1 => mux_o_831,
            S0 => ad(6)
        );

    mux_inst_861: MUX2
        port map (
            O => mux_o_861,
            I0 => mux_o_832,
            I1 => mux_o_833,
            S0 => ad(6)
        );

    mux_inst_862: MUX2
        port map (
            O => mux_o_862,
            I0 => mux_o_834,
            I1 => mux_o_835,
            S0 => ad(6)
        );

    mux_inst_863: MUX2
        port map (
            O => mux_o_863,
            I0 => mux_o_836,
            I1 => mux_o_837,
            S0 => ad(6)
        );

    mux_inst_864: MUX2
        port map (
            O => mux_o_864,
            I0 => mux_o_838,
            I1 => mux_o_839,
            S0 => ad(6)
        );

    mux_inst_865: MUX2
        port map (
            O => mux_o_865,
            I0 => mux_o_840,
            I1 => mux_o_841,
            S0 => ad(6)
        );

    mux_inst_866: MUX2
        port map (
            O => mux_o_866,
            I0 => mux_o_842,
            I1 => mux_o_843,
            S0 => ad(6)
        );

    mux_inst_867: MUX2
        port map (
            O => mux_o_867,
            I0 => mux_o_844,
            I1 => mux_o_845,
            S0 => ad(6)
        );

    mux_inst_868: MUX2
        port map (
            O => mux_o_868,
            I0 => mux_o_846,
            I1 => mux_o_847,
            S0 => ad(6)
        );

    mux_inst_869: MUX2
        port map (
            O => mux_o_869,
            I0 => mux_o_848,
            I1 => mux_o_849,
            S0 => ad(6)
        );

    mux_inst_870: MUX2
        port map (
            O => mux_o_870,
            I0 => mux_o_850,
            I1 => mux_o_851,
            S0 => ad(6)
        );

    mux_inst_871: MUX2
        port map (
            O => mux_o_871,
            I0 => mux_o_852,
            I1 => mux_o_853,
            S0 => ad(6)
        );

    mux_inst_872: MUX2
        port map (
            O => mux_o_872,
            I0 => mux_o_854,
            I1 => mux_o_855,
            S0 => ad(6)
        );

    mux_inst_873: MUX2
        port map (
            O => mux_o_873,
            I0 => mux_o_856,
            I1 => mux_o_857,
            S0 => ad(6)
        );

    mux_inst_874: MUX2
        port map (
            O => mux_o_874,
            I0 => mux_o_858,
            I1 => mux_o_859,
            S0 => ad(7)
        );

    mux_inst_875: MUX2
        port map (
            O => mux_o_875,
            I0 => mux_o_860,
            I1 => mux_o_861,
            S0 => ad(7)
        );

    mux_inst_876: MUX2
        port map (
            O => mux_o_876,
            I0 => mux_o_862,
            I1 => mux_o_863,
            S0 => ad(7)
        );

    mux_inst_877: MUX2
        port map (
            O => mux_o_877,
            I0 => mux_o_864,
            I1 => mux_o_865,
            S0 => ad(7)
        );

    mux_inst_878: MUX2
        port map (
            O => mux_o_878,
            I0 => mux_o_866,
            I1 => mux_o_867,
            S0 => ad(7)
        );

    mux_inst_879: MUX2
        port map (
            O => mux_o_879,
            I0 => mux_o_868,
            I1 => mux_o_869,
            S0 => ad(7)
        );

    mux_inst_880: MUX2
        port map (
            O => mux_o_880,
            I0 => mux_o_870,
            I1 => mux_o_871,
            S0 => ad(7)
        );

    mux_inst_881: MUX2
        port map (
            O => mux_o_881,
            I0 => mux_o_872,
            I1 => mux_o_873,
            S0 => ad(7)
        );

    mux_inst_882: MUX2
        port map (
            O => mux_o_882,
            I0 => mux_o_874,
            I1 => mux_o_875,
            S0 => ad(8)
        );

    mux_inst_883: MUX2
        port map (
            O => mux_o_883,
            I0 => mux_o_876,
            I1 => mux_o_877,
            S0 => ad(8)
        );

    mux_inst_884: MUX2
        port map (
            O => mux_o_884,
            I0 => mux_o_878,
            I1 => mux_o_879,
            S0 => ad(8)
        );

    mux_inst_885: MUX2
        port map (
            O => mux_o_885,
            I0 => mux_o_880,
            I1 => mux_o_881,
            S0 => ad(8)
        );

    mux_inst_886: MUX2
        port map (
            O => mux_o_886,
            I0 => mux_o_882,
            I1 => mux_o_883,
            S0 => ad(9)
        );

    mux_inst_887: MUX2
        port map (
            O => mux_o_887,
            I0 => mux_o_884,
            I1 => mux_o_885,
            S0 => ad(9)
        );

    mux_inst_888: MUX2
        port map (
            O => dout(6),
            I0 => mux_o_886,
            I1 => mux_o_887,
            S0 => ad(10)
        );

    mux_inst_889: MUX2
        port map (
            O => mux_o_889,
            I0 => ram16s_inst_1_dout(7),
            I1 => ram16s_inst_3_dout(7),
            S0 => ad(4)
        );

    mux_inst_890: MUX2
        port map (
            O => mux_o_890,
            I0 => ram16s_inst_5_dout(7),
            I1 => ram16s_inst_7_dout(7),
            S0 => ad(4)
        );

    mux_inst_891: MUX2
        port map (
            O => mux_o_891,
            I0 => ram16s_inst_9_dout(7),
            I1 => ram16s_inst_11_dout(7),
            S0 => ad(4)
        );

    mux_inst_892: MUX2
        port map (
            O => mux_o_892,
            I0 => ram16s_inst_13_dout(7),
            I1 => ram16s_inst_15_dout(7),
            S0 => ad(4)
        );

    mux_inst_893: MUX2
        port map (
            O => mux_o_893,
            I0 => ram16s_inst_17_dout(7),
            I1 => ram16s_inst_19_dout(7),
            S0 => ad(4)
        );

    mux_inst_894: MUX2
        port map (
            O => mux_o_894,
            I0 => ram16s_inst_21_dout(7),
            I1 => ram16s_inst_23_dout(7),
            S0 => ad(4)
        );

    mux_inst_895: MUX2
        port map (
            O => mux_o_895,
            I0 => ram16s_inst_25_dout(7),
            I1 => ram16s_inst_27_dout(7),
            S0 => ad(4)
        );

    mux_inst_896: MUX2
        port map (
            O => mux_o_896,
            I0 => ram16s_inst_29_dout(7),
            I1 => ram16s_inst_31_dout(7),
            S0 => ad(4)
        );

    mux_inst_897: MUX2
        port map (
            O => mux_o_897,
            I0 => ram16s_inst_33_dout(7),
            I1 => ram16s_inst_35_dout(7),
            S0 => ad(4)
        );

    mux_inst_898: MUX2
        port map (
            O => mux_o_898,
            I0 => ram16s_inst_37_dout(7),
            I1 => ram16s_inst_39_dout(7),
            S0 => ad(4)
        );

    mux_inst_899: MUX2
        port map (
            O => mux_o_899,
            I0 => ram16s_inst_41_dout(7),
            I1 => ram16s_inst_43_dout(7),
            S0 => ad(4)
        );

    mux_inst_900: MUX2
        port map (
            O => mux_o_900,
            I0 => ram16s_inst_45_dout(7),
            I1 => ram16s_inst_47_dout(7),
            S0 => ad(4)
        );

    mux_inst_901: MUX2
        port map (
            O => mux_o_901,
            I0 => ram16s_inst_49_dout(7),
            I1 => ram16s_inst_51_dout(7),
            S0 => ad(4)
        );

    mux_inst_902: MUX2
        port map (
            O => mux_o_902,
            I0 => ram16s_inst_53_dout(7),
            I1 => ram16s_inst_55_dout(7),
            S0 => ad(4)
        );

    mux_inst_903: MUX2
        port map (
            O => mux_o_903,
            I0 => ram16s_inst_57_dout(7),
            I1 => ram16s_inst_59_dout(7),
            S0 => ad(4)
        );

    mux_inst_904: MUX2
        port map (
            O => mux_o_904,
            I0 => ram16s_inst_61_dout(7),
            I1 => ram16s_inst_63_dout(7),
            S0 => ad(4)
        );

    mux_inst_905: MUX2
        port map (
            O => mux_o_905,
            I0 => ram16s_inst_65_dout(7),
            I1 => ram16s_inst_67_dout(7),
            S0 => ad(4)
        );

    mux_inst_906: MUX2
        port map (
            O => mux_o_906,
            I0 => ram16s_inst_69_dout(7),
            I1 => ram16s_inst_71_dout(7),
            S0 => ad(4)
        );

    mux_inst_907: MUX2
        port map (
            O => mux_o_907,
            I0 => ram16s_inst_73_dout(7),
            I1 => ram16s_inst_75_dout(7),
            S0 => ad(4)
        );

    mux_inst_908: MUX2
        port map (
            O => mux_o_908,
            I0 => ram16s_inst_77_dout(7),
            I1 => ram16s_inst_79_dout(7),
            S0 => ad(4)
        );

    mux_inst_909: MUX2
        port map (
            O => mux_o_909,
            I0 => ram16s_inst_81_dout(7),
            I1 => ram16s_inst_83_dout(7),
            S0 => ad(4)
        );

    mux_inst_910: MUX2
        port map (
            O => mux_o_910,
            I0 => ram16s_inst_85_dout(7),
            I1 => ram16s_inst_87_dout(7),
            S0 => ad(4)
        );

    mux_inst_911: MUX2
        port map (
            O => mux_o_911,
            I0 => ram16s_inst_89_dout(7),
            I1 => ram16s_inst_91_dout(7),
            S0 => ad(4)
        );

    mux_inst_912: MUX2
        port map (
            O => mux_o_912,
            I0 => ram16s_inst_93_dout(7),
            I1 => ram16s_inst_95_dout(7),
            S0 => ad(4)
        );

    mux_inst_913: MUX2
        port map (
            O => mux_o_913,
            I0 => ram16s_inst_97_dout(7),
            I1 => ram16s_inst_99_dout(7),
            S0 => ad(4)
        );

    mux_inst_914: MUX2
        port map (
            O => mux_o_914,
            I0 => ram16s_inst_101_dout(7),
            I1 => ram16s_inst_103_dout(7),
            S0 => ad(4)
        );

    mux_inst_915: MUX2
        port map (
            O => mux_o_915,
            I0 => ram16s_inst_105_dout(7),
            I1 => ram16s_inst_107_dout(7),
            S0 => ad(4)
        );

    mux_inst_916: MUX2
        port map (
            O => mux_o_916,
            I0 => ram16s_inst_109_dout(7),
            I1 => ram16s_inst_111_dout(7),
            S0 => ad(4)
        );

    mux_inst_917: MUX2
        port map (
            O => mux_o_917,
            I0 => ram16s_inst_113_dout(7),
            I1 => ram16s_inst_115_dout(7),
            S0 => ad(4)
        );

    mux_inst_918: MUX2
        port map (
            O => mux_o_918,
            I0 => ram16s_inst_117_dout(7),
            I1 => ram16s_inst_119_dout(7),
            S0 => ad(4)
        );

    mux_inst_919: MUX2
        port map (
            O => mux_o_919,
            I0 => ram16s_inst_121_dout(7),
            I1 => ram16s_inst_123_dout(7),
            S0 => ad(4)
        );

    mux_inst_920: MUX2
        port map (
            O => mux_o_920,
            I0 => ram16s_inst_125_dout(7),
            I1 => ram16s_inst_127_dout(7),
            S0 => ad(4)
        );

    mux_inst_921: MUX2
        port map (
            O => mux_o_921,
            I0 => ram16s_inst_129_dout(7),
            I1 => ram16s_inst_131_dout(7),
            S0 => ad(4)
        );

    mux_inst_922: MUX2
        port map (
            O => mux_o_922,
            I0 => ram16s_inst_133_dout(7),
            I1 => ram16s_inst_135_dout(7),
            S0 => ad(4)
        );

    mux_inst_923: MUX2
        port map (
            O => mux_o_923,
            I0 => ram16s_inst_137_dout(7),
            I1 => ram16s_inst_139_dout(7),
            S0 => ad(4)
        );

    mux_inst_924: MUX2
        port map (
            O => mux_o_924,
            I0 => ram16s_inst_141_dout(7),
            I1 => ram16s_inst_143_dout(7),
            S0 => ad(4)
        );

    mux_inst_925: MUX2
        port map (
            O => mux_o_925,
            I0 => ram16s_inst_145_dout(7),
            I1 => ram16s_inst_147_dout(7),
            S0 => ad(4)
        );

    mux_inst_926: MUX2
        port map (
            O => mux_o_926,
            I0 => ram16s_inst_149_dout(7),
            I1 => ram16s_inst_151_dout(7),
            S0 => ad(4)
        );

    mux_inst_927: MUX2
        port map (
            O => mux_o_927,
            I0 => ram16s_inst_153_dout(7),
            I1 => ram16s_inst_155_dout(7),
            S0 => ad(4)
        );

    mux_inst_928: MUX2
        port map (
            O => mux_o_928,
            I0 => ram16s_inst_157_dout(7),
            I1 => ram16s_inst_159_dout(7),
            S0 => ad(4)
        );

    mux_inst_929: MUX2
        port map (
            O => mux_o_929,
            I0 => ram16s_inst_161_dout(7),
            I1 => ram16s_inst_163_dout(7),
            S0 => ad(4)
        );

    mux_inst_930: MUX2
        port map (
            O => mux_o_930,
            I0 => ram16s_inst_165_dout(7),
            I1 => ram16s_inst_167_dout(7),
            S0 => ad(4)
        );

    mux_inst_931: MUX2
        port map (
            O => mux_o_931,
            I0 => ram16s_inst_169_dout(7),
            I1 => ram16s_inst_171_dout(7),
            S0 => ad(4)
        );

    mux_inst_932: MUX2
        port map (
            O => mux_o_932,
            I0 => ram16s_inst_173_dout(7),
            I1 => ram16s_inst_175_dout(7),
            S0 => ad(4)
        );

    mux_inst_933: MUX2
        port map (
            O => mux_o_933,
            I0 => ram16s_inst_177_dout(7),
            I1 => ram16s_inst_179_dout(7),
            S0 => ad(4)
        );

    mux_inst_934: MUX2
        port map (
            O => mux_o_934,
            I0 => ram16s_inst_181_dout(7),
            I1 => ram16s_inst_183_dout(7),
            S0 => ad(4)
        );

    mux_inst_935: MUX2
        port map (
            O => mux_o_935,
            I0 => ram16s_inst_185_dout(7),
            I1 => ram16s_inst_187_dout(7),
            S0 => ad(4)
        );

    mux_inst_936: MUX2
        port map (
            O => mux_o_936,
            I0 => ram16s_inst_189_dout(7),
            I1 => ram16s_inst_191_dout(7),
            S0 => ad(4)
        );

    mux_inst_937: MUX2
        port map (
            O => mux_o_937,
            I0 => ram16s_inst_193_dout(7),
            I1 => ram16s_inst_195_dout(7),
            S0 => ad(4)
        );

    mux_inst_938: MUX2
        port map (
            O => mux_o_938,
            I0 => ram16s_inst_197_dout(7),
            I1 => ram16s_inst_199_dout(7),
            S0 => ad(4)
        );

    mux_inst_939: MUX2
        port map (
            O => mux_o_939,
            I0 => ram16s_inst_201_dout(7),
            I1 => ram16s_inst_203_dout(7),
            S0 => ad(4)
        );

    mux_inst_940: MUX2
        port map (
            O => mux_o_940,
            I0 => ram16s_inst_205_dout(7),
            I1 => ram16s_inst_207_dout(7),
            S0 => ad(4)
        );

    mux_inst_941: MUX2
        port map (
            O => mux_o_941,
            I0 => ram16s_inst_209_dout(7),
            I1 => ram16s_inst_211_dout(7),
            S0 => ad(4)
        );

    mux_inst_942: MUX2
        port map (
            O => mux_o_942,
            I0 => ram16s_inst_213_dout(7),
            I1 => ram16s_inst_215_dout(7),
            S0 => ad(4)
        );

    mux_inst_943: MUX2
        port map (
            O => mux_o_943,
            I0 => ram16s_inst_217_dout(7),
            I1 => ram16s_inst_219_dout(7),
            S0 => ad(4)
        );

    mux_inst_944: MUX2
        port map (
            O => mux_o_944,
            I0 => ram16s_inst_221_dout(7),
            I1 => ram16s_inst_223_dout(7),
            S0 => ad(4)
        );

    mux_inst_945: MUX2
        port map (
            O => mux_o_945,
            I0 => ram16s_inst_225_dout(7),
            I1 => ram16s_inst_227_dout(7),
            S0 => ad(4)
        );

    mux_inst_946: MUX2
        port map (
            O => mux_o_946,
            I0 => ram16s_inst_229_dout(7),
            I1 => ram16s_inst_231_dout(7),
            S0 => ad(4)
        );

    mux_inst_947: MUX2
        port map (
            O => mux_o_947,
            I0 => ram16s_inst_233_dout(7),
            I1 => ram16s_inst_235_dout(7),
            S0 => ad(4)
        );

    mux_inst_948: MUX2
        port map (
            O => mux_o_948,
            I0 => ram16s_inst_237_dout(7),
            I1 => ram16s_inst_239_dout(7),
            S0 => ad(4)
        );

    mux_inst_949: MUX2
        port map (
            O => mux_o_949,
            I0 => ram16s_inst_241_dout(7),
            I1 => ram16s_inst_243_dout(7),
            S0 => ad(4)
        );

    mux_inst_950: MUX2
        port map (
            O => mux_o_950,
            I0 => ram16s_inst_245_dout(7),
            I1 => ram16s_inst_247_dout(7),
            S0 => ad(4)
        );

    mux_inst_951: MUX2
        port map (
            O => mux_o_951,
            I0 => ram16s_inst_249_dout(7),
            I1 => ram16s_inst_251_dout(7),
            S0 => ad(4)
        );

    mux_inst_952: MUX2
        port map (
            O => mux_o_952,
            I0 => ram16s_inst_253_dout(7),
            I1 => ram16s_inst_255_dout(7),
            S0 => ad(4)
        );

    mux_inst_953: MUX2
        port map (
            O => mux_o_953,
            I0 => mux_o_889,
            I1 => mux_o_890,
            S0 => ad(5)
        );

    mux_inst_954: MUX2
        port map (
            O => mux_o_954,
            I0 => mux_o_891,
            I1 => mux_o_892,
            S0 => ad(5)
        );

    mux_inst_955: MUX2
        port map (
            O => mux_o_955,
            I0 => mux_o_893,
            I1 => mux_o_894,
            S0 => ad(5)
        );

    mux_inst_956: MUX2
        port map (
            O => mux_o_956,
            I0 => mux_o_895,
            I1 => mux_o_896,
            S0 => ad(5)
        );

    mux_inst_957: MUX2
        port map (
            O => mux_o_957,
            I0 => mux_o_897,
            I1 => mux_o_898,
            S0 => ad(5)
        );

    mux_inst_958: MUX2
        port map (
            O => mux_o_958,
            I0 => mux_o_899,
            I1 => mux_o_900,
            S0 => ad(5)
        );

    mux_inst_959: MUX2
        port map (
            O => mux_o_959,
            I0 => mux_o_901,
            I1 => mux_o_902,
            S0 => ad(5)
        );

    mux_inst_960: MUX2
        port map (
            O => mux_o_960,
            I0 => mux_o_903,
            I1 => mux_o_904,
            S0 => ad(5)
        );

    mux_inst_961: MUX2
        port map (
            O => mux_o_961,
            I0 => mux_o_905,
            I1 => mux_o_906,
            S0 => ad(5)
        );

    mux_inst_962: MUX2
        port map (
            O => mux_o_962,
            I0 => mux_o_907,
            I1 => mux_o_908,
            S0 => ad(5)
        );

    mux_inst_963: MUX2
        port map (
            O => mux_o_963,
            I0 => mux_o_909,
            I1 => mux_o_910,
            S0 => ad(5)
        );

    mux_inst_964: MUX2
        port map (
            O => mux_o_964,
            I0 => mux_o_911,
            I1 => mux_o_912,
            S0 => ad(5)
        );

    mux_inst_965: MUX2
        port map (
            O => mux_o_965,
            I0 => mux_o_913,
            I1 => mux_o_914,
            S0 => ad(5)
        );

    mux_inst_966: MUX2
        port map (
            O => mux_o_966,
            I0 => mux_o_915,
            I1 => mux_o_916,
            S0 => ad(5)
        );

    mux_inst_967: MUX2
        port map (
            O => mux_o_967,
            I0 => mux_o_917,
            I1 => mux_o_918,
            S0 => ad(5)
        );

    mux_inst_968: MUX2
        port map (
            O => mux_o_968,
            I0 => mux_o_919,
            I1 => mux_o_920,
            S0 => ad(5)
        );

    mux_inst_969: MUX2
        port map (
            O => mux_o_969,
            I0 => mux_o_921,
            I1 => mux_o_922,
            S0 => ad(5)
        );

    mux_inst_970: MUX2
        port map (
            O => mux_o_970,
            I0 => mux_o_923,
            I1 => mux_o_924,
            S0 => ad(5)
        );

    mux_inst_971: MUX2
        port map (
            O => mux_o_971,
            I0 => mux_o_925,
            I1 => mux_o_926,
            S0 => ad(5)
        );

    mux_inst_972: MUX2
        port map (
            O => mux_o_972,
            I0 => mux_o_927,
            I1 => mux_o_928,
            S0 => ad(5)
        );

    mux_inst_973: MUX2
        port map (
            O => mux_o_973,
            I0 => mux_o_929,
            I1 => mux_o_930,
            S0 => ad(5)
        );

    mux_inst_974: MUX2
        port map (
            O => mux_o_974,
            I0 => mux_o_931,
            I1 => mux_o_932,
            S0 => ad(5)
        );

    mux_inst_975: MUX2
        port map (
            O => mux_o_975,
            I0 => mux_o_933,
            I1 => mux_o_934,
            S0 => ad(5)
        );

    mux_inst_976: MUX2
        port map (
            O => mux_o_976,
            I0 => mux_o_935,
            I1 => mux_o_936,
            S0 => ad(5)
        );

    mux_inst_977: MUX2
        port map (
            O => mux_o_977,
            I0 => mux_o_937,
            I1 => mux_o_938,
            S0 => ad(5)
        );

    mux_inst_978: MUX2
        port map (
            O => mux_o_978,
            I0 => mux_o_939,
            I1 => mux_o_940,
            S0 => ad(5)
        );

    mux_inst_979: MUX2
        port map (
            O => mux_o_979,
            I0 => mux_o_941,
            I1 => mux_o_942,
            S0 => ad(5)
        );

    mux_inst_980: MUX2
        port map (
            O => mux_o_980,
            I0 => mux_o_943,
            I1 => mux_o_944,
            S0 => ad(5)
        );

    mux_inst_981: MUX2
        port map (
            O => mux_o_981,
            I0 => mux_o_945,
            I1 => mux_o_946,
            S0 => ad(5)
        );

    mux_inst_982: MUX2
        port map (
            O => mux_o_982,
            I0 => mux_o_947,
            I1 => mux_o_948,
            S0 => ad(5)
        );

    mux_inst_983: MUX2
        port map (
            O => mux_o_983,
            I0 => mux_o_949,
            I1 => mux_o_950,
            S0 => ad(5)
        );

    mux_inst_984: MUX2
        port map (
            O => mux_o_984,
            I0 => mux_o_951,
            I1 => mux_o_952,
            S0 => ad(5)
        );

    mux_inst_985: MUX2
        port map (
            O => mux_o_985,
            I0 => mux_o_953,
            I1 => mux_o_954,
            S0 => ad(6)
        );

    mux_inst_986: MUX2
        port map (
            O => mux_o_986,
            I0 => mux_o_955,
            I1 => mux_o_956,
            S0 => ad(6)
        );

    mux_inst_987: MUX2
        port map (
            O => mux_o_987,
            I0 => mux_o_957,
            I1 => mux_o_958,
            S0 => ad(6)
        );

    mux_inst_988: MUX2
        port map (
            O => mux_o_988,
            I0 => mux_o_959,
            I1 => mux_o_960,
            S0 => ad(6)
        );

    mux_inst_989: MUX2
        port map (
            O => mux_o_989,
            I0 => mux_o_961,
            I1 => mux_o_962,
            S0 => ad(6)
        );

    mux_inst_990: MUX2
        port map (
            O => mux_o_990,
            I0 => mux_o_963,
            I1 => mux_o_964,
            S0 => ad(6)
        );

    mux_inst_991: MUX2
        port map (
            O => mux_o_991,
            I0 => mux_o_965,
            I1 => mux_o_966,
            S0 => ad(6)
        );

    mux_inst_992: MUX2
        port map (
            O => mux_o_992,
            I0 => mux_o_967,
            I1 => mux_o_968,
            S0 => ad(6)
        );

    mux_inst_993: MUX2
        port map (
            O => mux_o_993,
            I0 => mux_o_969,
            I1 => mux_o_970,
            S0 => ad(6)
        );

    mux_inst_994: MUX2
        port map (
            O => mux_o_994,
            I0 => mux_o_971,
            I1 => mux_o_972,
            S0 => ad(6)
        );

    mux_inst_995: MUX2
        port map (
            O => mux_o_995,
            I0 => mux_o_973,
            I1 => mux_o_974,
            S0 => ad(6)
        );

    mux_inst_996: MUX2
        port map (
            O => mux_o_996,
            I0 => mux_o_975,
            I1 => mux_o_976,
            S0 => ad(6)
        );

    mux_inst_997: MUX2
        port map (
            O => mux_o_997,
            I0 => mux_o_977,
            I1 => mux_o_978,
            S0 => ad(6)
        );

    mux_inst_998: MUX2
        port map (
            O => mux_o_998,
            I0 => mux_o_979,
            I1 => mux_o_980,
            S0 => ad(6)
        );

    mux_inst_999: MUX2
        port map (
            O => mux_o_999,
            I0 => mux_o_981,
            I1 => mux_o_982,
            S0 => ad(6)
        );

    mux_inst_1000: MUX2
        port map (
            O => mux_o_1000,
            I0 => mux_o_983,
            I1 => mux_o_984,
            S0 => ad(6)
        );

    mux_inst_1001: MUX2
        port map (
            O => mux_o_1001,
            I0 => mux_o_985,
            I1 => mux_o_986,
            S0 => ad(7)
        );

    mux_inst_1002: MUX2
        port map (
            O => mux_o_1002,
            I0 => mux_o_987,
            I1 => mux_o_988,
            S0 => ad(7)
        );

    mux_inst_1003: MUX2
        port map (
            O => mux_o_1003,
            I0 => mux_o_989,
            I1 => mux_o_990,
            S0 => ad(7)
        );

    mux_inst_1004: MUX2
        port map (
            O => mux_o_1004,
            I0 => mux_o_991,
            I1 => mux_o_992,
            S0 => ad(7)
        );

    mux_inst_1005: MUX2
        port map (
            O => mux_o_1005,
            I0 => mux_o_993,
            I1 => mux_o_994,
            S0 => ad(7)
        );

    mux_inst_1006: MUX2
        port map (
            O => mux_o_1006,
            I0 => mux_o_995,
            I1 => mux_o_996,
            S0 => ad(7)
        );

    mux_inst_1007: MUX2
        port map (
            O => mux_o_1007,
            I0 => mux_o_997,
            I1 => mux_o_998,
            S0 => ad(7)
        );

    mux_inst_1008: MUX2
        port map (
            O => mux_o_1008,
            I0 => mux_o_999,
            I1 => mux_o_1000,
            S0 => ad(7)
        );

    mux_inst_1009: MUX2
        port map (
            O => mux_o_1009,
            I0 => mux_o_1001,
            I1 => mux_o_1002,
            S0 => ad(8)
        );

    mux_inst_1010: MUX2
        port map (
            O => mux_o_1010,
            I0 => mux_o_1003,
            I1 => mux_o_1004,
            S0 => ad(8)
        );

    mux_inst_1011: MUX2
        port map (
            O => mux_o_1011,
            I0 => mux_o_1005,
            I1 => mux_o_1006,
            S0 => ad(8)
        );

    mux_inst_1012: MUX2
        port map (
            O => mux_o_1012,
            I0 => mux_o_1007,
            I1 => mux_o_1008,
            S0 => ad(8)
        );

    mux_inst_1013: MUX2
        port map (
            O => mux_o_1013,
            I0 => mux_o_1009,
            I1 => mux_o_1010,
            S0 => ad(9)
        );

    mux_inst_1014: MUX2
        port map (
            O => mux_o_1014,
            I0 => mux_o_1011,
            I1 => mux_o_1012,
            S0 => ad(9)
        );

    mux_inst_1015: MUX2
        port map (
            O => dout(7),
            I0 => mux_o_1013,
            I1 => mux_o_1014,
            S0 => ad(10)
        );

end Behavioral; --Gowin_RAM16S
